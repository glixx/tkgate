//: version "2.1-a2"
//: property prefix = "_GG"

//: /netlistBegin main
module main;    //: root_module
reg w6;    //: /sn:0 {0}(98,88)(114,88)(114,88)(131,88){1}
reg w7;    //: /sn:0 {0}(101,243)(117,243)(117,243)(134,243){1}
reg w16;    //: /sn:0 {0}(451,75)(467,75)(467,75)(484,75){1}
reg w14;    //: /sn:0 {0}(97,377)(138,377)(138,406){1}
reg w19;    //: /sn:0 {0}(484,141)(468,141)(468,141)(451,141){1}
reg w15;    //: /sn:0 {0}(451,109)(492,109)(492,136){1}
reg w4;    //: /sn:0 {0}(101,209)(142,209)(142,238){1}
reg w3;    //: /sn:0 {0}(101,277)(142,277)(142,304){1}
reg w21;    //: /sn:0 {0}(453,234)(469,234)(469,234)(486,234){1}
reg w24;    //: /sn:0 {0}(453,268)(494,268)(494,295){1}
reg w23;    //: /sn:0 {0}(486,300)(470,300)(470,300)(453,300){1}
reg w1;    //: /sn:0 {0}(98,54)(139,54)(139,83){1}
reg w22;    //: /sn:0 {0}(453,200)(494,200)(494,229){1}
reg w17;    //: /sn:0 {0}(451,41)(492,41)(492,70){1}
reg w12;    //: /sn:0 {0}(130,477)(114,477)(114,477)(97,477){1}
reg w2;    //: /sn:0 {0}(98,122)(139,122)(139,149){1}
reg w10;    //: /sn:0 {0}(97,445)(138,445)(138,472){1}
reg w13;    //: /sn:0 {0}(97,411)(113,411)(113,411)(130,411){1}
reg w5;    //: /sn:0 /dp:1 {0}(131,154)(115,154)(115,154)(98,154){1}
reg w9;    //: /sn:0 {0}(134,309)(118,309)(118,309)(101,309){1}
wire w0;    //: /sn:0 {0}(147,88)(162,88)(162,121){1}
//: {2}(164,123)(194,123)(194,107){3}
//: {4}(162,125)(162,154)(147,154){5}
tri1 w20;    //: /sn:0 /dp:3 {0}(502,234)(517,234)(517,267){1}
//: {2}(519,269)(570,269)(570,249){3}
//: {4}(517,271)(517,300)(502,300){5}
tri0 w18;    //: /sn:0 /dp:3 {0}(500,75)(515,75)(515,108){1}
//: {2}(517,110)(566,110)(566,90){3}
//: {4}(515,112)(515,141)(500,141){5}
wand w8;    //: /sn:0 /dp:3 {0}(150,243)(165,243)(165,276){1}
//: {2}(167,278)(193,278)(193,268){3}
//: {4}(165,280)(165,309)(150,309){5}
wor w11;    //: /sn:0 /dp:3 {0}(146,411)(161,411)(161,444){1}
//: {2}(163,446)(191,446)(191,424){3}
//: {4}(161,448)(161,477)(146,477){5}
//: enddecls

  //: SWITCH g8 (w3) @(84,277) /sn:0 /w:[ 0 ] /st:0
  //: SWITCH g4 (w2) @(81,122) /sn:0 /w:[ 0 ] /st:0
  //: SWITCH g37 (w24) @(436,268) /sn:0 /w:[ 0 ] /st:0
  _GGBUFIF #(4, 6) g34 (.Z(w20), .I(w23), .E(w24));   //: @(492,300) /sn:0 /w:[ 5 0 1 ]
  //: joint g13 (w8) @(165, 278) /w:[ 2 1 -1 4 ]
  //: SWITCH g3 (w1) @(81,54) /sn:0 /w:[ 0 ] /st:0
  //: SWITCH g2 (w6) @(81,88) /sn:0 /w:[ 0 ] /st:0
  _GGBUFIF #(4, 6) g1 (.Z(w0), .I(w5), .E(w2));   //: @(137,154) /sn:0 /w:[ 5 0 1 ]
  //: SWITCH g16 (w10) @(80,445) /sn:0 /w:[ 0 ] /st:0
  _GGBUFIF #(4, 6) g11 (.Z(w8), .I(w9), .E(w3));   //: @(140,309) /sn:0 /w:[ 5 0 1 ]
  _GGBUFIF #(4, 6) g28 (.Z(w18), .I(w16), .E(w17));   //: @(490,75) /sn:0 /w:[ 0 1 1 ]
  //: SWITCH g10 (w7) @(84,243) /sn:0 /w:[ 0 ] /st:0
  _GGBUFIF #(4, 6) g32 (.Z(w20), .I(w21), .E(w22));   //: @(492,234) /sn:0 /w:[ 0 1 1 ]
  //: joint g27 (w18) @(515, 110) /w:[ 2 1 -1 4 ]
  //: SWITCH g19 (w13) @(80,411) /sn:0 /w:[ 0 ] /st:0
  //: SWITCH g38 (w22) @(436,200) /sn:0 /w:[ 0 ] /st:0
  //: LED g6 (w0) @(194,100) /sn:0 /w:[ 3 ] /type:0
  //: SWITCH g9 (w4) @(84,209) /sn:0 /w:[ 0 ] /st:0
  //: joint g7 (w0) @(162, 123) /w:[ 2 1 -1 4 ]
  _GGBUFIF #(4, 6) g31 (.Z(w18), .I(w19), .E(w15));   //: @(490,141) /sn:0 /w:[ 5 0 1 ]
  //: SWITCH g20 (w14) @(80,377) /sn:0 /w:[ 0 ] /st:0
  _GGBUFIF #(4, 6) g15 (.Z(w8), .I(w7), .E(w4));   //: @(140,243) /sn:0 /w:[ 0 1 1 ]
  //: SWITCH g39 (w23) @(436,300) /sn:0 /w:[ 1 ] /st:0
  //: LED g29 (w18) @(566,83) /sn:0 /w:[ 3 ] /type:0
  //: SWITCH g25 (w16) @(434,75) /sn:0 /w:[ 0 ] /st:0
  //: joint g17 (w11) @(161, 446) /w:[ 2 1 -1 4 ]
  //: SWITCH g14 (w9) @(84,309) /sn:0 /w:[ 1 ] /st:0
  //: SWITCH g5 (w5) @(81,154) /sn:0 /w:[ 1 ] /st:0
  //: LED g36 (w20) @(570,242) /sn:0 /w:[ 3 ] /type:0
  //: SWITCH g24 (w15) @(434,109) /sn:0 /w:[ 0 ] /st:0
  _GGBUFIF #(4, 6) g21 (.Z(w11), .I(w13), .E(w14));   //: @(136,411) /sn:0 /w:[ 0 1 1 ]
  //: LED g23 (w11) @(191,417) /sn:0 /w:[ 3 ] /type:0
  //: SWITCH g35 (w21) @(436,234) /sn:0 /w:[ 0 ] /st:0
  //: SWITCH g26 (w17) @(434,41) /sn:0 /w:[ 0 ] /st:0
  //: SWITCH g22 (w12) @(80,477) /sn:0 /w:[ 1 ] /st:0
  _GGBUFIF #(4, 6) g0 (.Z(w0), .I(w6), .E(w1));   //: @(137,88) /sn:0 /w:[ 0 1 1 ]
  _GGBUFIF #(4, 6) g18 (.Z(w11), .I(w12), .E(w10));   //: @(136,477) /sn:0 /w:[ 5 0 1 ]
  //: LED g12 (w8) @(193,261) /sn:0 /w:[ 3 ] /type:0
  //: joint g33 (w20) @(517, 269) /w:[ 2 1 -1 4 ]
  //: SWITCH g30 (w19) @(434,141) /sn:0 /w:[ 1 ] /st:0

endmodule
//: /netlistEnd

//: /builtinBegin
module _GGBUFIF #(.Dez(1), .Diz(1)) (Z, I, E);
input E;
input I;
output Z;

  specify
    (E *> Z) = Dez;
    (I *> Z) = Diz;
  endspecify

  assign Z = E ? (I) : 1'bz;

endmodule
//: /builtinEnd

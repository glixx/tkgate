//: version "2.1-a2"
//: property prefix = "_GG"
//: property title = "module_tut.v"

//: /netlistBegin main
module main;    //: root_module
//: enddecls

  //: comment g0 @(23,20) /sn:0
  //: /line:"<h3 color=blue>Creating a Module Definition</h3>"
  //: /line:""
  //: /line:"1) Press <img src=\"blk_new.gif\"> on the tool bar."
  //: /line:""
  //: /line:"2) Enter the name of the new module."
  //: /line:""
  //: /line:"3) Select the type of module (Netlist or HDL)"
  //: /line:""
  //: /line:"4) Click \"OK\" to create the module."
  //: /line:""
  //: /line:"5) Edit it by double clicking on it in the module list."
  //: /line:""
  //: /line:"<a href=\"module_tut.v\">Click here to return to the main module tutorial.</a>"
  //: /end

endmodule
//: /netlistEnd

//: version "2.1-a2"
//: property prefix = "_GG"
//: property title = "module_tut.v"

//: /netlistBegin main
module main;    //: root_module
//: enddecls

  //: comment g0 @(23,20) /sn:0
  //: /line:"<h3 color=blue>Erzeugen einer Moduldefinition</h3>"
  //: /line:""
  //: /line:"1) Drücke <img src=\"blk_new.gif\"> auf der Toolbar."
  //: /line:""
  //: /line:"2) Gib den Namen des neuen Moduls ein."
  //: /line:""
  //: /line:"3) Wähle den Modultyp (Netzliste oder HDL)"
  //: /line:""
  //: /line:"4) Klicke \"OK\" und erzeuge das Modul."
  //: /line:""
  //: /line:"5) Editiere esdurch Doppelklick in der Modulliste."
  //: /line:""
  //: /line:"<a href=\"module_tut.v\">Hier klicken, um ins Hauptmenu zurückzukehren.</a>"
  //: /end

endmodule
//: /netlistEnd

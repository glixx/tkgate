//: version "2.1-a2"
//: property encoding = "utf-8"
//: property locale = "ru"
//: property prefix = "_GG"
//: property title = "index.v"
//: property showSwitchNets = 0
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
//: enddecls

  //: comment g4 @(553,317) /sn:0 /anc:1
  //: /line:"<h3><a href=\"ex6/coke.v\"><img src=example_coke.gif>"
  //: /line:"Автомат газировки</a></h3>"
  //: /line:"Этот пример использует механизм"
  //: /line:"виртуальных периферийных устройств (ВПУ)"
  //: /line:"TkGate для создания интерактивной модели"
  //: /line:"\"Автомат газировки\", которой можно управлять"
  //: /line:"с помощью пользовательской схемы."
  //: /line:"Включена только модель. Сможете ли Вы построить"
  //: /line:"контроллер для неё?"
  //: /line:""
  //: /end
  //: comment g3 @(32,317) /sn:0 /anc:1
  //: /line:"<a href=\"ex4/trff.v\"><img src=\"example_trff.gif\">"
  //: /line:"<h3>Защёлка на уровне транзисторов</h3></a>"
  //: /line:"Триггер, реализованный с"
  //: /line:"использованием Н-МОП и П-МОП"
  //: /line:"элементов."
  //: /line:""
  //: /end
  //: comment g2 @(551,30) /sn:0 /anc:1
  //: /line:"<a href=\"ex3/counter.v\"><img src=\"example_counter.gif\">"
  //: /line:"<h3>8-разрядный счётчик</h3></a>"
  //: /line:"Счётчик, реализованный с"
  //: /line:"использованием регистра и"
  //: /line:"сумматора."
  //: /end
  //: comment g1 @(299,30) /sn:0 /anc:1
  //: /line:"<a href=\"ex2/flipflop.v\"><img src=\"example_flipflop.gif\">"
  //: /line:"<h3>4-разрядный счётчик</h3></a>"
  //: /line:"4-разрядный счётчик, реализованный с"
  //: /line:"использованием четырёх одноразрядных"
  //: /line:"D-защёлок."
  //: /end
  //: comment g6 @(20,552) /sn:0
  //: /line:"<font size=5><a href=\"@T/welcome.v\">Вернуться на главную страницу</a></font>"
  //: /end
  //: comment g7 @(787,27) /sn:0
  //: /line:"<a href=\"ex7/stdlogic.v\"><img src=\"example_counter.gif\">"
  //: /line:"<h3>Микросхемы 74xx</h3></a>"
  //: /line:"Несколько примеров схем с"
  //: /line:"использованием библиотеки"
  //: /line:"микросхем стандартной логики"
  //: /line:"серии 74."
  //: /end
  //: comment g5 @(301,317) /sn:0 /anc:1
  //: /line:"<h3><a href=\"ex5/menagerie.v\"><img src=\"example_menagerie.gif\">"
  //: /line:"Компьютер \"Зверинец\"</a></h3>"
  //: /line:"Простой микропроцессор с микрокодом,"
  //: /line:"который выполняет игру \"Животные\""
  //: /line:"во время симуляции."
  //: /end
  //: comment g0 @(32,30) /sn:0 /anc:1
  //: /line:"<h3><a href=\"ex1/combinational.v\"><img src=\"example_combinational.gif\">"
  //: /line:"Комбинационная логика</a></h3>"
  //: /line:"Простой 3-разрядный сумматор, который"
  //: /line:"можно запускать в симуляторе."
  //: /line:"Нажмите кнопку запуска, затем"
  //: /line:"изменяйте значения переключателей и"
  //: /line:"смотрите, как меняются состояния"
  //: /line:"светодиодов."
  //: /line:""
  //: /end

endmodule
//: /netlistEnd


`timescale 1ns/1ns


//: version "2.0-b10"
//: property encoding = "iso8859-1"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "stdlogic.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"
//: require "74xx"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg [15:0] A_NET;    //: {0}(#:-101,129)(#:50:-173,129){1}
reg w3;    //: /sn:0 {0}(314,199)(227,199)(227,192)(33,192)(33,366){1}
//: {2}(35,368)(51,368){3}
//: {4}(53,366)(53,199)(119,199){5}
//: {6}(53,370)(53,563)(119,563){7}
//: {8}(31,368)(-190,368){9}
//: {10}(33,370)(33,559)(354,559){11}
reg [3:0] w18;    //: /sn:0 {0}(#:-139,290)(#:-172,290){1}
supply0 w2;    //: /sn:0 {0}(62,163)(62,183)(119,183){1}
wire w6;    //: /sn:0 {0}(119,167)(104,167){1}
wire w32;    //: /sn:0 {0}(-95,164)(-3,164)(-3,467)(119,467){1}
wire w7;    //: /sn:0 {0}(119,151)(104,151){1}
wire w45;    //: /sn:0 {0}(354,607)(264,607)(264,392)(167,392)(167,331){1}
//: {2}(169,329)(260,329)(260,247)(314,247){3}
//: {4}(165,329)(48,329)(48,297){5}
//: {6}(48,293)(48,247)(119,247){7}
//: {8}(46,295)(-74,295){9}
//: {10}(-78,295)(-133,295){11}
//: {12}(-76,297)(-76,611)(119,611){13}
wire w73;    //: /sn:0 {0}(354,511)(334,511){1}
wire w93;    //: /sn:0 {0}(409,87)(523,87)(523,240)(599,240){1}
wire w96;    //: /sn:0 {0}(214,435)(238,435)(238,377)(482,377)(482,270)(599,270){1}
wire w46;    //: /sn:0 {0}(314,231)(251,231)(251,319)(203,319){1}
//: {2}(199,319)(39,319)(39,287){3}
//: {4}(39,283)(39,231)(119,231){5}
//: {6}(37,285)(-64,285){7}
//: {8}(-68,285)(-133,285){9}
//: {10}(-66,287)(-66,595)(119,595){11}
//: {12}(201,321)(201,381)(272,381)(272,591)(354,591){13}
wire w60;    //: /sn:0 {0}(119,547)(89,547)(89,359)(446,359)(446,135)(409,135){1}
wire w61;    //: /sn:0 {0}(409,119)(424,119){1}
wire w99;    //: /sn:0 {0}(599,300)(515,300)(515,415)(449,415){1}
wire w14;    //: /sn:0 {0}(214,167)(229,167){1}
wire w16;    //: /sn:0 {0}(214,135)(252,135)(252,183)(314,183){1}
wire w56;    //: /sn:0 {0}(-95,104)(-54,104)(-54,-49)(285,-49)(285,71)(314,71){1}
wire w15;    //: /sn:0 {0}(214,151)(229,151){1}
wire w19;    //: /sn:0 {0}(214,87)(248,87)(248,23)(563,23)(563,200)(599,200){1}
wire w81;    //: /sn:0 {0}(449,511)(464,511){1}
wire w38;    //: /sn:0 {0}(214,499)(299,499)(299,543)(354,543){1}
wire w51;    //: /sn:0 {0}(314,151)(299,151){1}
wire w0;    //: /sn:0 {0}(354,623)(236,623)(236,399)(148,399)(148,340){1}
//: {2}(150,338)(271,338)(271,263)(314,263){3}
//: {4}(146,338)(57,338)(57,307){5}
//: {6}(57,303)(57,263)(119,263){7}
//: {8}(55,305)(-89,305){9}
//: {10}(-93,305)(-133,305){11}
//: {12}(-91,307)(-91,627)(119,627){13}
wire w97;    //: /sn:0 {0}(214,451)(249,451)(249,388)(492,388)(492,280)(599,280){1}
wire w37;    //: /sn:0 {0}(214,515)(229,515){1}
wire w64;    //: /sn:0 {0}(409,71)(534,71)(534,230)(599,230){1}
wire w34;    //: /sn:0 {0}(-95,144)(12,144)(12,435)(119,435){1}
wire w21;    //: /sn:0 {0}(214,55)(226,55)(226,-1)(584,-1)(584,180)(599,180){1}
wire w43;    //: /sn:0 {0}(214,419)(229,419)(229,368)(473,368)(473,260)(599,260){1}
wire w75;    //: /sn:0 {0}(354,479)(339,479){1}
wire w76;    //: /sn:0 {0}(354,463)(331,463)(331,694)(-36,694)(-36,204)(-95,204){1}
wire w102;    //: /sn:0 {0}(449,463)(550,463)(550,330)(599,330){1}
wire w54;    //: /sn:0 {0}(-95,124)(-30,124)(-30,-25)(265,-25)(265,103)(314,103){1}
wire w31;    //: /sn:0 {0}(119,483)(104,483){1}
wire w58;    //: /sn:0 {0}(409,167)(424,167){1}
wire w90;    //: /sn:0 {0}(214,103)(259,103)(259,33)(552,33)(552,210)(599,210){1}
wire w100;    //: /sn:0 {0}(449,431)(526,431)(526,310)(599,310){1}
wire w28;    //: /sn:0 {0}(119,531)(104,531){1}
wire w20;    //: /sn:0 {0}(214,71)(237,71)(237,12)(574,12)(574,190)(599,190){1}
wire w36;    //: /sn:0 {0}(214,531)(229,531){1}
wire w1;    //: /sn:0 {0}(354,575)(282,575)(282,353)(229,353)(229,313){1}
//: {2}(231,311)(246,311)(246,215)(314,215){3}
//: {4}(227,311)(29,311)(29,277){5}
//: {6}(29,273)(29,215)(119,215){7}
//: {8}(27,275)(-55,275){9}
//: {10}(-59,275)(-133,275){11}
//: {12}(-57,277)(-57,579)(119,579){13}
wire w82;    //: /sn:0 {0}(632,467)(632,495)(449,495){1}
wire w65;    //: /sn:0 {0}(409,55)(543,55)(543,220)(599,220){1}
wire w74;    //: /sn:0 {0}(354,495)(339,495){1}
wire w98;    //: /sn:0 {0}(599,290)(502,290)(502,397)(259,397)(259,467)(214,467){1}
wire w8;    //: /sn:0 {0}(119,135)(104,135){1}
wire w35;    //: /sn:0 {0}(-95,134)(22,134)(22,419)(119,419){1}
wire w30;    //: /sn:0 {0}(119,499)(104,499){1}
wire w101;    //: /sn:0 {0}(599,320)(536,320)(536,447)(449,447){1}
wire w17;    //: /sn:0 {0}(214,119)(229,119){1}
wire w53;    //: /sn:0 {0}(314,119)(299,119){1}
wire w59;    //: /sn:0 {0}(409,151)(424,151){1}
wire w62;    //: /sn:0 {0}(409,103)(514,103)(514,250)(599,250){1}
wire w11;    //: /sn:0 {0}(-95,74)(94,74)(94,87)(119,87){1}
wire w12;    //: /sn:0 {0}(-95,64)(104,64)(104,71)(119,71){1}
wire w57;    //: /sn:0 {0}(-95,94)(-66,94)(-66,-61)(295,-61)(295,55)(314,55){1}
wire w77;    //: /sn:0 {0}(354,447)(321,447)(321,685)(-25,685)(-25,194)(-95,194){1}
wire w83;    //: /sn:0 {0}(449,479)(464,479){1}
wire w10;    //: /sn:0 {0}(-95,84)(87,84)(87,103)(119,103){1}
wire w78;    //: /sn:0 {0}(-95,184)(-17,184)(-17,676)(313,676)(313,431)(354,431){1}
wire w13;    //: /sn:0 {0}(-95,54)(104,54)(104,55)(119,55){1}
wire w72;    //: /sn:0 {0}(354,527)(339,527){1}
wire [15:0] w27;    //: /sn:0 {0}(#:605,255)(640,255){1}
wire w33;    //: /sn:0 {0}(-95,154)(4,154)(4,451)(119,451){1}
wire w52;    //: /sn:0 {0}(314,135)(299,135){1}
wire w29;    //: /sn:0 {0}(119,515)(104,515){1}
wire w80;    //: /sn:0 {0}(449,527)(503,527){1}
wire w9;    //: /sn:0 {0}(119,119)(104,119){1}
wire w50;    //: /sn:0 {0}(314,167)(299,167){1}
wire w79;    //: /sn:0 {0}(-95,174)(-9,174)(-9,668)(304,668)(304,415)(354,415){1}
wire w39;    //: /sn:0 {0}(214,483)(229,483){1}
wire w55;    //: /sn:0 {0}(-95,114)(-42,114)(-42,-37)(275,-37)(275,87)(314,87){1}
//: enddecls

  //: joint g8 (w1) @(-57, 275) /w:[ 9 -1 10 12 ]
  //: LED g4 (w27) @(647,255) /sn:0 /R:3 /w:[ 1 ] /type:2
  //: joint g13 (w46) @(39, 285) /w:[ -1 4 6 3 ]
  H74181 g3 (._A0(w79), ._A1(w78), ._A2(w77), ._A3(w76), ._B0(w75), ._B1(w74), ._B2(w73), ._B3(w72), .Cn(w38), .M(w3), .S0(w1), .S1(w46), .S2(w45), .S3(w0), ._F0(w99), ._F1(w100), ._F2(w101), ._F3(w102), .AEB(w83), .CnP4(w82), ._G(w81), ._P(w80));   //: @(355, 399) /sz:(93, 240) /sn:0 /p:[ Li0>1 Li1>1 Li2>0 Li3>0 Li4>0 Li5>0 Li6>0 Li7>0 Li8>1 Li9>11 Li10>0 Li11>13 Li12>0 Li13>0 Ro0<1 Ro1<0 Ro2<1 Ro3<0 Ro4<0 Ro5<1 Ro6<0 Ro7<0 ]
  H74181 g2 (._A0(w57), ._A1(w56), ._A2(w55), ._A3(w54), ._B0(w53), ._B1(w52), ._B2(w51), ._B3(w50), .Cn(w16), .M(w3), .S0(w1), .S1(w46), .S2(w45), .S3(w0), ._F0(w65), ._F1(w64), ._F2(w93), ._F3(w62), .AEB(w61), .CnP4(w60), ._G(w59), ._P(w58));   //: @(315, 39) /sz:(93, 240) /sn:0 /p:[ Li0>1 Li1>1 Li2>1 Li3>1 Li4>0 Li5>0 Li6>0 Li7>0 Li8>1 Li9>0 Li10>3 Li11>0 Li12>3 Li13>3 Ro0<0 Ro1<0 Ro2<0 Ro3<0 Ro4<0 Ro5<1 Ro6<0 Ro7<0 ]
  H74181 g1 (._A0(w35), ._A1(w34), ._A2(w33), ._A3(w32), ._B0(w31), ._B1(w30), ._B2(w29), ._B3(w28), .Cn(w60), .M(w3), .S0(w1), .S1(w46), .S2(w45), .S3(w0), ._F0(w43), ._F1(w96), ._F2(w97), ._F3(w98), .AEB(w39), .CnP4(w38), ._G(w37), ._P(w36));   //: @(120, 403) /sz:(93, 240) /sn:0 /p:[ Li0>1 Li1>1 Li2>1 Li3>1 Li4>0 Li5>0 Li6>0 Li7>0 Li8>0 Li9>7 Li10>13 Li11>11 Li12>13 Li13>13 Ro0<0 Ro1<0 Ro2<0 Ro3<1 Ro4<0 Ro5<0 Ro6<0 Ro7<0 ]
  //: joint g16 (w1) @(229, 311) /w:[ 2 -1 4 1 ]
  //: joint g11 (w0) @(-91, 305) /w:[ 9 -1 10 12 ]
  //: DIP A (A_NET) @(-211,129) /R:1 /w:[ 1 ] /st:2 /dn:1
  //: joint g10 (w45) @(-76, 295) /w:[ 9 -1 10 12 ]
  //: joint g19 (w0) @(148, 338) /w:[ 2 -1 4 1 ]
  assign {w0, w45, w46, w1} = w18; //: CONCAT g6  @(-138,290) /sn:0 /R:2 /w:[ 11 11 9 11 0 ] /dr:0 /tp:1 /drp:0
  //: DIP OP (w18) @(-210,290) /R:1 /w:[ 1 ] /st:0 /dn:1
  //: joint g9 (w46) @(-66, 285) /w:[ 7 -1 8 10 ]
  assign {w76, w77, w78, w79, w32, w33, w34, w35, w54, w55, w56, w57, w10, w11, w12, w13} = A_NET; //: CONCAT g7  @(-100,129) /sn:0 /R:2 /w:[ 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 ] /dr:0 /tp:1 /drp:0
  //: GROUND g20 (w2) @(62,157) /sn:0 /R:2 /w:[ 0 ]
  //: joint g15 (w0) @(57, 305) /w:[ -1 6 8 5 ]
  //: joint g17 (w46) @(201, 319) /w:[ 1 -1 2 12 ]
  //: joint g14 (w45) @(48, 295) /w:[ -1 6 8 5 ]
  assign w27 = {w102, w101, w100, w99, w98, w97, w96, w43, w62, w93, w64, w65, w90, w19, w20, w21}; //: CONCAT g5  @(604,255) /sn:0 /w:[ 0 1 0 1 0 0 1 1 1 1 1 1 1 1 1 1 1 ] /dr:1 /tp:1 /drp:1
  //: joint g24 (w3) @(33, 368) /w:[ 2 1 8 10 ]
  //: LED g21 (w82) @(632,460) /sn:0 /w:[ 0 ] /type:0
  //: joint g23 (w3) @(53, 368) /w:[ -1 4 3 6 ]
  //: SWITCH g22 (w3) @(-207,368) /sn:0 /w:[ 9 ] /st:1 /dn:1
  H74181 g0 (._A0(w13), ._A1(w12), ._A2(w11), ._A3(w10), ._B0(w9), ._B1(w8), ._B2(w7), ._B3(w6), .Cn(w2), .M(w3), .S0(w1), .S1(w46), .S2(w45), .S3(w0), ._F0(w21), ._F1(w20), ._F2(w19), ._F3(w90), .AEB(w17), .CnP4(w16), ._G(w15), ._P(w14));   //: @(120, 39) /sz:(93, 240) /sn:0 /p:[ Li0>1 Li1>1 Li2>1 Li3>1 Li4>0 Li5>0 Li6>0 Li7>0 Li8>1 Li9>5 Li10>7 Li11>5 Li12>7 Li13>7 Ro0<0 Ro1<0 Ro2<0 Ro3<0 Ro4<0 Ro5<0 Ro6<0 Ro7<0 ]
  //: joint g18 (w45) @(167, 329) /w:[ 2 -1 4 1 ]
  //: joint g12 (w1) @(29, 275) /w:[ -1 6 8 5 ]

endmodule
//: /netlistEnd


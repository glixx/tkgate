//: version "2.1-a2"
//: property encoding = "utf-8"
//: property locale = "de"
//: property prefix = "_GG"
//: property title = "Tutorial page"
//: property showSwitchNets = 0
//: property discardChanges = 1
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin PAGE1
module PAGE1;    //: root_module
//: enddecls

  //: comment g1 @(475,291) /sn:0 /R:14 /anc:1
  //: /line:"<a href=\"welcome.v\">Zurück zur Hauptseite von TkGate.</a>"
  //: /end
  //: comment g0 @(476,49) /sn:0 /anc:1
  //: /line:"<a href=\"welcome.v\"><img src=\"biggatelogo.gif\"></a>"
  //: /end
  //: comment g18 @(10,10) /sn:0 /anc:1
  //: /line:"<h1>Lernabschnitte:</h1>"
  //: /line:""
  //: /line:"<h3><a href=\"create.v\">1. Erzeugen einer Schaltung</a></h3>"
  //: /line:""
  //: /line:"<h3><a href=\"gates.v\">2. Gatter editieren</a></h3> - Grundlagen zum Konfigurieren von Gattern."
  //: /line:""
  //: /line:"<h3><a href=\"wires.v\">3. Leitungen editieren</a></h3> - Grundlagen zum Konfigurieren von Leitungen."
  //: /line:""
  //: /line:"<h3><a href=\"group.v\">4. Editieren von Gattergruppen</a></h3>"
  //: /line:" - Bearbeiten von Gruppen benachbarter Gatter."
  //: /line:""
  //: /line:"<h3><a href=\"modules.v\">5. Benutzung von Modulen</a></h3>"
  //: /line:" - Verwenden von Modulkapselung in der Schaltung."
  //: /line:""
  //: /line:"<h3><a href=\"advanced.v\">6. Fortgeschrittene Editiertechniken</a></h3>"
  //: /line:" - Einige weniger gebräuchliche Editiertricks."
  //: /line:""
  //: /line:"<h3><a href=\"combinational1.v\">7. Simulation von Schaltnetzen</a></h3>"
  //: /line:" - Simulieren eines Schaltnetzes."
  //: /line:""
  //: /line:"<h3><a href=\"sequential1.v\">8. Simulation von Schaltwerken</a></h3> - Simulation sequentieller Schaltungen."
  //: /line:""
  //: /line:"<h3><a href=\"verilog.v\">9. Schaltungen mit Verilog-Text</a></h3> - Erzeugen von Modulen, die textuelle Verilog-Beschreibungen enthalten."
  //: /line:""
  //: /line:"<h3><a href=\"options.v\">10. Anpassen von TkGate</a></h3> - Konfigurieren nach eigenem Geschmack."
  //: /line:""
  //: /end

endmodule
//: /netlistEnd


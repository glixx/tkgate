//: version "2.1"
//: property prefix = "_GG"
//: property title = "greek.v"

//: /netlistBegin main
module main;    //: root_module
//: enddecls

  //: comment g1 @(195,37) /sn:0
  //: /line:"&alpha; alpha "
  //: /line:"&beta; beta "
  //: /line:"&gamma; gamma "
  //: /line:"&delta; delta "
  //: /line:"&epsilon; epsilon "
  //: /line:"&zeta; zeta "
  //: /line:"&eta; eta "
  //: /line:"&theta; theta "
  //: /line:"&iota; iota "
  //: /line:"&kappa; kappa "
  //: /line:"&lambda; lambda "
  //: /line:"&mu; mu "
  //: /line:"&nu; nu "
  //: /line:"&xi; xi "
  //: /line:"&omicron; omicron "
  //: /line:"&pi; pi "
  //: /line:"&rho; rho "
  //: /line:"&sigmaf; sigmaf "
  //: /line:"&sigma; sigma "
  //: /line:"&tau; tau "
  //: /line:"&upsilon; upsilon "
  //: /line:"&phi; phi "
  //: /line:"&chi; chi "
  //: /line:"&psi; psi "
  //: /line:"&omega; omega "
  //: /line:"&thetasym; thetasym "
  //: /line:"&upsih; upsih "
  //: /line:"&piv; piv  "
  //: /line:""
  //: /end
  //: comment g0 @(61,55) /sn:0
  //: /line:"&Alpha; Alpha "
  //: /line:"&Beta; Beta "
  //: /line:"&Gamma; Gamma "
  //: /line:"&Delta; Delta "
  //: /line:"&Epsilon; Epsilon "
  //: /line:"&Zeta; Zeta "
  //: /line:"&Eta; Eta "
  //: /line:"&Theta; Theta "
  //: /line:"&Iota; Iota "
  //: /line:"&Kappa; Kappa "
  //: /line:"&Lambda; Lambda "
  //: /line:"&Mu; Mu "
  //: /line:"&Nu; Nu "
  //: /line:"&Xi; Xi "
  //: /line:"&Omicron; Omicron "
  //: /line:"&Pi; Pi "
  //: /line:"&Rho; Rho "
  //: /line:"&Sigma; Sigma "
  //: /line:"&Tau; Tau "
  //: /line:"&Upsilon; Upsilon "
  //: /line:"&Phi; Phi "
  //: /line:"&Chi; Chi "
  //: /line:"&Psi; Psi "
  //: /line:"&Omega; Omega "
  //: /line:""
  //: /end

endmodule
//: /netlistEnd

//: version "2.1-a2"
//: property encoding = "utf-8"
//: property locale = "ru"
//: property prefix = "_GG"
//: property title = "Страница Учебного руководства"
//: property showSwitchNets = 0
//: property discardChanges = 1
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin PAGE1
module PAGE1;    //: root_module
//: enddecls

  //: comment g1 @(475,291) /sn:0 /R:14 /anc:1
  //: /line:"<a href=\"welcome.v\">Вернуться к стартовой схеме TkGate.</a>"
  //: /end
  //: comment g0 @(476,49) /sn:0 /anc:1
  //: /line:"<a href=\"welcome.v\"><img src=\"biggatelogo.gif\"></a>"
  //: /end
  //: comment g18 @(10,10) /sn:0 /anc:1
  //: /line:"<h1>Разделы руководства:</h1>"
  //: /line:""
  //: /line:"<h3><a href=\"create.v\">1. Создание схемы</a></h3> - Начните с создания простой схемы."
  //: /line:""
  //: /line:"<h3><a href=\"gates.v\">2. Редактирование вентилей</a></h3> - Основы редактирования вентилей."
  //: /line:""
  //: /line:"<h3><a href=\"wires.v\">3. Редактирование проводов</a></h3> - Основы редактирования проводов."
  //: /line:""
  //: /line:"<h3><a href=\"group.v\">4. Средства редактирования групп</a></h3> - Управляйте группами вентилей."
  //: /line:""
  //: /line:"<h3><a href=\"modules.v\">5. Использование модулей</a></h3> - Использование моделей в ваших схемах."
  //: /line:""
  //: /line:"<h3><a href=\"advanced.v\">6. Расширенные техники редактирования</a></h3> - Изучите особенности"
  //: /line:"и тонкости редактирования схем."
  //: /line:""
  //: /line:"<h3><a href=\"combinational1.v\">7. Комбинационная симуляция</a></h3> - Имитируйте работу схемы"
  //: /line:"с комбинационной логикой."
  //: /line:""
  //: /line:"<h3><a href=\"sequential1.v\">8. Последовательная симуляция</a></h3> - Имитируйте работу схемы с"
  //: /line:"последовательной логикой."
  //: /line:""
  //: /line:"<h3><a href=\"verilog.v\">9. Текстовый Verilog</a></h3> - Создавайте модули с текстовым описанием"
  //: /line:"на Verilog."
  //: /line:""
  //: /line:"<h3><a href=\"options.v\">10. Настройка TkGate</a></h3> - Настраивайте TkGate по своему вкусу."
  //: /line:""
  //: /end

endmodule
//: /netlistEnd


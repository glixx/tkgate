//: version "2.1-a2"
//: property prefix = "_GG"
//: property title = "sim_tut.v"
//: property useExtBars = 0
//: property discardChanges = 1

//: /netlistBegin main
module main;    //: root_module
//: enddecls

  //: frame g15 @(600,25) /sn:0 /wi:213 /ht:149 /tx:"Tutorials"
  //: comment g14 @(629,42) /sn:0
  //: /line:"<a href=\"welcome_tut.v\">TkGate Introduction</a><br>"
  //: /line:"<a href=\"create_tut.v\">Creating a Circuit</a><br>"
  //: /line:"<a href=\"edit1_tut.v\">Basic Editing Modes</a><br>"
  //: /line:"<a href=\"edit2_tut.v\">Group Editing Features</a><br>"
  //: /line:"<a href=\"edwire_tut.v\">Editing Wires</a><br>"
  //: /line:"<a href=\"module_tut.v\">Using Modules</a><br>"
  //: /line:"<a href=\"sim_tut.v\">Combinational Simulation</a><br>"
  //: /line:"<a href=\"seqsim_tut.v\">Sequential Simulation</a>"
  //: /end
  //: comment g0 @(21,26) /sn:0
  //: /line:"<h2>Glossary</h2>"
  //: /line:""
  //: /line:"<b>epoch</b>: The smallest unit of time understood by the simulator."
  //: /line:""
  //: /line:"<a name=verconst></a><b>Verilog format constant</b>: The first number indicates the bit width, the"
  //: /line:"letter indicates the radix, and the last number the value.  For example, the \"1\""
  //: /line:"in \"1'b0\" indicates that this is a 1-bit value, the \"b\" indicates the value is"
  //: /line:"given in binary, and the \"0\" indicates the value of the signal."
  //: /end

endmodule
//: /netlistEnd

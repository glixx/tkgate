//: version "2.2"
//: property encoding = "utf-8"
//: property locale = "ja"
//: property prefix = "_GG"
//: property title = "Tutorial page"
//: property showSwitchNets = 0
//: property discardChanges = 1
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin PAGE1
module PAGE1;    //: root_module
//: enddecls

  //: comment g1 @(475,291) /sn:0 /R:14 /anc:1
  //: /line:"<a href=\"welcome.v\">Go back to the TkGate main page.</a>"
  //: /end
  //: comment g0 @(476,49) /sn:0 /anc:1
  //: /line:"<a href=\"welcome.v\"><img src=\"biggatelogo.gif\"></a>"
  //: /end
  //: comment g18 @(10,10) /sn:0 /anc:1
  //: /line:"<font color=chocolate>Tutorial Chapters:</font>"
  //: /line:""
  //: /line:"<font color=purple><a href=\"create.v\">1. 回路の作成</a></font> - Get started by creating a simple circuit."
  //: /line:""
  //: /line:"<font color=purple><a href=\"gates.v\">2. Editing Gates</a></font> - The basics of editing gates."
  //: /line:""
  //: /line:"<font color=purple><a href=\"wires.v\">3. ワイヤの編集</a></font> - The basics of editing wires."
  //: /line:""
  //: /line:"<font color=purple><a href=\"group.v\">4. グループの編集機能</a></font> - Operate on groups of gates."
  //: /line:""
  //: /line:"<font color=purple><a href=\"modules.v\">5. モジュールの使い方</a></font> - Using modules in your circuit."
  //: /line:""
  //: /line:"<font color=purple><a href=\"advanced.v\">6. Advanced Editing Techniques</a></font> - Learn advanced editing tricks."
  //: /line:""
  //: /line:"<font color=purple><a href=\"combinational1.v\">7. 組合せ回路のシミュレーション</a></font> - Simulate a circuit with"
  //: /line:"combinational logic."
  //: /line:""
  //: /line:"<font color=purple><a href=\"sequential1.v\">8. 順序回路のシミュレーション</a></font> - Simulate a circuit with sequential logic."
  //: /line:""
  //: /line:"<font color=purple><a href=\"verilog.v\">9. Textual Verilog</a></font> - Create modules with textual Verilog descriptions."
  //: /line:""
  //: /line:"<font color=purple><a href=\"options.v\">10. Customizing TkGate</a></font> - Customize TkGate to suit your tastes."
  //: /line:""
  //: /end

endmodule
//: /netlistEnd


//: version "2.1"
//: property encoding = "utf-8"
//: property locale = "de"
//: property prefix = "_GG"
//: property title = "Customizing TkGate"
//: property showSwitchNets = 0
//: property discardChanges = 1
//: property timingViolationMode = 2
//: property initTime = "0 ns"
//: require "tty"

`timescale 1ns/1ns

//: /netlistBegin PAGE1
module PAGE1;    //: root_module
//: enddecls

  //: comment g1 @(219,134) /sn:0 /anc:1
  //: /line:"<img src=iface.gif>"
  //: /end
  //: comment g9 @(10,10) /anc:1
  //: /line:"<h3>Anpassen von TkGate</h3>"
  //: /line:""
  //: /line:"Dieser Abschnitt führt einige der Optionen ein, mit denen TkGate angepaßt werden kann."
  //: /line:"Die Definitionen der Optionen werden in einer Datei namens \".tkgate2-preferences\" im"
  //: /line:"Heimatverzeichnis gespeichert."
  //: /end
  //: comment g0 @(10,310) /sn:0 /anc:1
  //: /line:"<tutorial-navigation>"
  //: /end

endmodule
//: /netlistEnd

//: /netlistBegin PAGE3
module PAGE3();
//: interface  /sz:(40, 40) /bd:[ ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
//: enddecls

  //: comment g1 @(134,181) /sn:0 /anc:1
  //: /line:"<img src=example_bindings.gif>"
  //: /end
  //: comment g9 @(10,10) /anc:1
  //: /line:"<h3>Anpassen von TkGate</h3> <b>(Setzen der Tastaturbindungen)</b>"
  //: /line:""
  //: /line:"Man kann die Tastaturbindungen für die Benutzung der <font color=red2>Schnittstelle</font> Taste der Optionen-Dialogbox"
  //: /line:"anpassen. Zur Zeit kann man zwischen \"emacs\"-style und \"Windows\"-Stil wählen. Das paßt"
  //: /line:"die Tastaturbelegungen für Operationen wie Ausschneiden/Einfügen an die Gepflogenheiten von emacs oder Windows an."
  //: /line:"Die Tastenbelegungen für die Erzeugung von Gattern bleiben allerdings erhalten."
  //: /end
  //: comment g0 @(10,310) /sn:0
  //: /line:"<tutorial-navigation>"
  //: /end

endmodule
//: /netlistEnd

//: /netlistBegin PAGE2
module PAGE2();
//: interface  /sz:(40, 40) /bd:[ ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
//: enddecls

  //: comment g1 @(116,149) /sn:0 /anc:1
  //: /line:"<img src=example_name.gif>"
  //: /end
  //: comment g9 @(10,10) /anc:1
  //: /line:"<h3>Anpassen von TkGate</h3> <b>(Angabe der persönlichen Daten)</b>"
  //: /line:""
  //: /line:"Zum Festlegen der TkGate Optionen öffnet man die Optionen Dialogbox durch Auswahl von <font color=red2>Datei &rarr; Optionen</font> aus dem"
  //: /line:"Hauptmenu. Gib den Namen der Institution und den Benutzernamen in der \"Organisation\" Dialogbox ein. Die eingegebenen Werte"
  //: /line:"werden in jeder Druckausgabe von TkGate-Schaltungen benutzt."
  //: /end
  //: comment g0 @(10,310) /sn:0 /anc:1
  //: /line:"<tutorial-navigation>"
  //: /end

endmodule
//: /netlistEnd


//: version "2.1"
//: property encoding = "utf-8"
//: property locale = "uk"
//: property prefix = "_GG"
//: property title = "Example page"
//: property showSwitchNets = 0
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
//: enddecls

  //: comment g4 @(553,317) /sn:0 /anc:1
  //: /line:"<a href=\"ex6/coke.v\"><img src=example_coke.gif>"
  //: /line:"<h3>Coke Machine</h3></a>"
  //: /line:"This example uses TkGate's Viritual"
  //: /line:"Peripheral Device (VPD) mechanism to"
  //: /line:"create an interactive \"Coke Machine\""
  //: /line:"that can be controlled by a user circuit."
  //: /line:"Only the coke machine device itself is"
  //: /line:"included. Can you build a controller"
  //: /line:"for it?"
  //: /line:""
  //: /end
  //: comment g3 @(32,317) /sn:0 /anc:1
  //: /line:"<a href=\"ex4/trff.v\"><img src=\"example_trff.gif\">"
  //: /line:"<h3>Transistor-Level FF</h3></a>"
  //: /line:"A flop-flop implemented using"
  //: /line:"nmos and pmos devices."
  //: /line:""
  //: /end
  //: comment g2 @(551,30) /sn:0 /anc:1
  //: /line:"<a href=\"ex3/counter.v\"><img src=\"example_counter.gif\">"
  //: /line:"<h3>8-бітовий лічильник</h3></a>"
  //: /line:"A counter implemented using the"
  //: /line:"register and adder devices."
  //: /end
  //: comment g1 @(299,30) /sn:0 /anc:1
  //: /line:"<a href=\"ex2/flipflop.v\"><img src=\"example_flipflop.gif\">"
  //: /line:"<h3>4-бітовий лічильник</h3></a>"
  //: /line:"A 4-bitcounter implemented using"
  //: /line:"four single-bit D-flip-flops."
  //: /end
  //: comment g6 @(20,552) /sn:0
  //: /line:"<font size=5><a href=\"@T/welcome.v\">Go back to the TkGate main page</a></font>"
  //: /end
  //: comment g7 @(787,27) /sn:0
  //: /line:"<a href=\"ex7/stdlogic.v\"><img src=\"example_counter.gif\">"
  //: /line:"<h3>Microcircuits 74xx</h3></a>"
  //: /line:"A few examples of circuits"
  //: /line:"using the standard"
  //: /line:"74 series"
  //: /line:"logic circuit library."
  //: /end
  //: comment g5 @(301,317) /sn:0 /anc:1
  //: /line:"<a href=\"ex5/menagerie.v\"><img src=\"example_menagerie.gif\">"
  //: /line:"<h3>Menagerie CPU</h3></a>"
  //: /line:"A simple microcode-based CPU that"
  //: /line:"will play the \"Animals\" game on a"
  //: /line:"TTY device when simulated."
  //: /end
  //: comment g0 @(32,30) /sn:0 /anc:1
  //: /line:"<a href=\"ex1/combinational.v\"><img src=\"example_combinational.gif\">"
  //: /line:"<h3>Combinational Logic</h3></a>"
  //: /line:"A simple 3-bit adder that you"
  //: /line:"simulate. Push the play button"
  //: /line:"then click on the switches and"
  //: /line:"watch how the LEDs change."
  //: /line:""
  //: /end

endmodule
//: /netlistEnd


`timescale 1ns/1ns


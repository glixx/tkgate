//: version "2.0-b10"
//: property encoding = "utf-8"
//: property locale = "ru"
//: property prefix = "_GG"
//: property title = "stdlogic.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"
//: require "74xx"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg [15:0] A_NET;    //: {0}(#:50:62,167)(192,167){1}
//: {2}(196,167)(249,167){3}
//: {4}(#:194,169)(194,346)(243,346){5}
reg w0;    //: /sn:0 {0}(17,373)(128,373){1}
//: {2}(130,371)(130,215)(249,215){3}
//: {4}(130,375)(130,394)(243,394){5}
reg w3;    //: /sn:0 {0}(19,316)(142,316){1}
//: {2}(144,314)(144,199)(249,199){3}
//: {4}(144,318)(144,378)(243,378){5}
reg [3:0] w18;    //: /sn:0 {0}(#:45,410)(93,410){1}
//: {2}(97,410)(243,410){3}
//: {4}(95,408)(95,231)(249,231){5}
reg [15:0] w2;    //: /sn:0 {0}(#:61,221)(85,221)(85,183)(157,183){1}
//: {2}(161,183)(50:249,183){3}
//: {4}(#:159,185)(159,362)(243,362){5}
wire [15:0] w4;    //: /sn:0 {0}(#:449,183)(393,183){1}
wire w11;    //: /sn:0 {0}(475,318)(475,346)(441,346){1}
wire [15:0] w10;    //: /sn:0 {0}(#:490,362)(441,362){1}
wire w5;    //: /sn:0 {0}(393,167)(433,167)(433,129){1}
//: enddecls

  //: SWITCH M (w0) @(0,373) /w:[ 0 ] /st:0 /dn:1
  //: joint g4 (A_NET) @(194, 167) /w:[ 2 -1 1 4 ]
  //: joint g8 (w0) @(130, 373) /w:[ -1 2 1 4 ]
  ALU16_74181_74182 g3 (.A(A_NET), .B(w2), .CI(w3), .M(w0), .OP(w18), .CO(w11), .F(w10));   //: @(244, 330) /sz:(196, 96) /sn:0 /p:[ Li0>5 Li1>5 Li2>5 Li3>5 Li4>3 Ro0<1 Ro1<1 ]
  //: comment g2 @(58,18) /sn:0
  //: /line:"00 - НЕ <b>A</b>"
  //: /line:"05 - НЕ <b>B</b>"
  //: /line:"06 - <b>A</b> ИСКЛ. ИЛИ <b>B</b>"
  //: /line:"0B - <b>A</b> И <b>B</b>"
  //: /line:"0С - <b>A</b> ИЛИ <b>B</b>"
  //: /end
  //: LED g1 (w5) @(433,122) /sn:0 /w:[ 1 ] /type:0
  //: DIP B_DIP (w2) @(23,221) /R:1 /w:[ 0 ] /st:244 /dn:1
  //: DIP OP_DIP (w18) @(7,410) /R:1 /w:[ 0 ] /st:9 /dn:1
  //: LED g11 (w10) @(497,362) /sn:0 /R:3 /w:[ 0 ] /type:2
  //: LED g10 (w11) @(475,311) /sn:0 /w:[ 0 ] /type:0
  //: LED g6 (w4) @(456,183) /sn:0 /R:3 /w:[ 0 ] /type:2
  //: joint g7 (w3) @(144, 316) /w:[ -1 2 1 4 ]
  //: joint g9 (w18) @(95, 410) /w:[ 2 4 1 -1 ]
  //: SWITCH CI (w3) @(2,316) /w:[ 0 ] /st:1 /dn:1
  //: joint g5 (w2) @(159, 183) /w:[ 2 -1 1 4 ]
  ALU16_74181 g0 (.A(A_NET), .B(w2), .CI(w3), .M(w0), .S(w18), .CO(w5), .F(w4));   //: @(250, 151) /sz:(142, 96) /sn:0 /p:[ Li0>3 Li1>3 Li2>3 Li3>3 Li4>5 Ro0<0 Ro1<1 ]
  //: DIP A_DIP (A_NET) @(24,167) /R:1 /w:[ 0 ] /st:171 /dn:1

endmodule
//: /netlistEnd

//: /netlistBegin ALU16_74181
module ALU16_74181(F, S, M, B, CI, CO, A);
//: interface  /sz:(142, 96) /bd:[ Li0>A[15:0](16/96) Li1>B[15:0](32/96) Li2>CI(48/96) Li3>M(64/96) Li4>S[3:0](80/96) Ro0<CO(16/96) Ro1<F[15:0](32/96) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input M;    //: {0}(519,556)(353,556)(353,695)(19,695)(19,565){1}
//: {2}(21,563)(71,563)(71,563)(120,563){3}
//: {4}(19,561)(19,465)(18,465)(18,370){5}
//: {6}(18,366)(18,327){7}
//: {8}(20,325)(429,325)(429,189)(519,189){9}
//: {10}(18,323)(18,189)(120,189){11}
//: {12}(16,368)(-194,368)(-194,368)(99:-406,368){13}
input [15:0] B;    //: /sn:0 {0}(#:-331,559)(#:-406,559){1}
output [15:0] F;    //: /sn:0 {0}(1048,256)(#:986,256){1}
input [15:0] A;    //: {0}(#:80:-406,79)(-373,79)(-373,79)(#:58:-331,79){1}
output CO;    //: /sn:0 {0}(1025,491)(819,491)(819,492)(614,492){1}
input CI;    //: /sn:0 {0}(120,173)(-347,173)(-347,218)(-406,218){1}
input [3:0] S;    //: {0}(#:70:-406,290)(-367,290)(-367,290)(#:-331,290){1}
wire w32;    //: /sn:0 {0}(-325,114)(-249,114)(-249,467)(120,467){1}
wire w6;    //: /sn:0 {0}(120,157)(-171,157)(-171,514)(-325,514){1}
wire w73;    //: /sn:0 {0}(519,508)(386,508)(386,789)(-169,789)(-169,624)(-325,624){1}
wire w45;    //: /sn:0 {0}(519,604)(471,604)(471,355)(216,355)(216,297){1}
//: {2}(218,295)(466,295)(466,237)(519,237){3}
//: {4}(214,295)(50,295){5}
//: {6}(48,293)(48,237)(120,237){7}
//: {8}(46,295)(-15,295){9}
//: {10}(-19,295)(-325,295){11}
//: {12}(-17,297)(-17,611)(120,611){13}
wire w93;    //: /sn:0 {0}(614,77)(906,77)(906,241)(980,241){1}
wire w96;    //: /sn:0 {0}(215,435)(288,435)(288,736)(863,736)(863,271)(980,271){1}
wire w7;    //: /sn:0 {0}(120,141)(-182,141)(-182,504)(-325,504){1}
wire w46;    //: /sn:0 {0}(519,221)(453,221)(453,285)(227,285){1}
//: {2}(223,285)(41,285){3}
//: {4}(39,283)(39,221)(120,221){5}
//: {6}(37,285)(-4,285){7}
//: {8}(-8,285)(-325,285){9}
//: {10}(-6,287)(-6,595)(120,595){11}
//: {12}(225,287)(225,346)(481,346)(481,588)(519,588){13}
wire w99;    //: /sn:0 {0}(980,301)(893,301)(893,412)(614,412){1}
wire w61;    //: /sn:0 {0}(614,109)(629,109){1}
wire w60;    //: /sn:0 {0}(120,547)(35,547)(35,706)(841,706)(841,125)(614,125){1}
wire w56;    //: /sn:0 {0}(-325,54)(-170,54)(-170,-109)(397,-109)(397,61)(519,61){1}
wire w16;    //: /sn:0 {0}(215,125)(310,125)(310,173)(519,173){1}
wire w14;    //: /sn:0 {0}(215,157)(230,157){1}
wire w81;    //: /sn:0 {0}(614,508)(629,508){1}
wire w19;    //: /sn:0 {0}(215,77)(297,77)(297,6)(945,6)(945,201)(980,201){1}
wire w15;    //: /sn:0 {0}(215,141)(230,141){1}
wire w38;    //: /sn:0 {0}(215,499)(251,499)(251,540)(519,540){1}
wire w51;    //: /sn:0 {0}(-325,544)(-104,544)(-104,-46)(336,-46)(336,141)(519,141){1}
wire w0;    //: /sn:0 {0}(519,620)(460,620)(460,363)(207,363)(207,307){1}
//: {2}(209,305)(478,305)(478,253)(519,253){3}
//: {4}(205,305)(59,305){5}
//: {6}(57,303)(57,253)(120,253){7}
//: {8}(55,305)(-25,305){9}
//: {10}(-29,305)(-325,305){11}
//: {12}(-27,307)(-27,627)(120,627){13}
wire w97;    //: /sn:0 {0}(215,451)(277,451)(277,747)(875,747)(875,281)(980,281){1}
wire w64;    //: /sn:0 {0}(614,61)(917,61)(917,231)(980,231){1}
wire w37;    //: /sn:0 {0}(215,515)(230,515){1}
wire w34;    //: /sn:0 {0}(-325,94)(-227,94)(-227,435)(120,435){1}
wire w76;    //: /sn:0 {0}(519,460)(343,460)(343,683)(-288,683)(-288,154)(-325,154){1}
wire w75;    //: /sn:0 {0}(519,476)(363,476)(363,765)(-148,765)(-148,604)(-325,604){1}
wire w102;    //: /sn:0 {0}(614,460)(922,460)(922,331)(980,331){1}
wire w43;    //: /sn:0 {0}(215,419)(299,419)(299,726)(851,726)(851,261)(980,261){1}
wire w21;    //: /sn:0 {0}(215,45)(273,45)(273,-19)(966,-19)(966,181)(980,181){1}
wire w54;    //: /sn:0 {0}(-325,74)(-144,74)(-144,-85)(370,-85)(370,93)(519,93){1}
wire w100;    //: /sn:0 {0}(614,428)(902,428)(902,311)(980,311){1}
wire w58;    //: /sn:0 {0}(614,157)(629,157){1}
wire w31;    //: /sn:0 {0}(-325,564)(-77,564)(-77,483)(120,483){1}
wire w90;    //: /sn:0 {0}(215,93)(308,93)(308,21)(934,21)(934,211)(980,211){1}
wire w28;    //: /sn:0 {0}(120,531)(-39,531)(-39,594)(-325,594){1}
wire w36;    //: /sn:0 {0}(215,531)(230,531){1}
wire w20;    //: /sn:0 {0}(215,61)(285,61)(285,-6)(956,-6)(956,191)(980,191){1}
wire w1;    //: /sn:0 {0}(519,572)(490,572)(490,336)(233,336)(233,277){1}
//: {2}(235,275)(441,275)(441,205)(519,205){3}
//: {4}(231,275)(31,275){5}
//: {6}(29,273)(29,205)(120,205){7}
//: {8}(27,275)(6,275){9}
//: {10}(2,275)(-325,275){11}
//: {12}(4,277)(4,579)(120,579){13}
wire w74;    //: /sn:0 {0}(519,492)(374,492)(374,776)(-159,776)(-159,614)(-325,614){1}
wire w65;    //: /sn:0 {0}(614,45)(926,45)(926,221)(980,221){1}
wire w98;    //: /sn:0 {0}(980,291)(887,291)(887,756)(264,756)(264,467)(215,467){1}
wire w40;    //: /sn:0 {0}(120,515)(-50,515)(-50,584)(-325,584){1}
wire w35;    //: /sn:0 {0}(-325,84)(-215,84)(-215,419)(120,419){1}
wire w8;    //: /sn:0 {0}(120,125)(-195,125)(-195,494)(-325,494){1}
wire w101;    //: /sn:0 {0}(980,321)(912,321)(912,444)(614,444){1}
wire w30;    //: /sn:0 {0}(120,499)(-64,499)(-64,574)(-325,574){1}
wire w17;    //: /sn:0 {0}(215,109)(230,109){1}
wire w53;    //: /sn:0 {0}(519,109)(358,109)(358,-72)(-130,-72)(-130,524)(-325,524){1}
wire w59;    //: /sn:0 {0}(614,141)(629,141){1}
wire w62;    //: /sn:0 {0}(614,93)(897,93)(897,251)(980,251){1}
wire w57;    //: /sn:0 {0}(-325,44)(-182,44)(-182,-121)(409,-121)(409,45)(519,45){1}
wire w12;    //: /sn:0 {0}(-325,14)(94,14)(94,61)(120,61){1}
wire w11;    //: /sn:0 {0}(-325,24)(80,24)(80,77)(120,77){1}
wire w77;    //: /sn:0 {0}(519,444)(333,444)(333,672)(-279,672)(-279,144)(-325,144){1}
wire w83;    //: /sn:0 {0}(614,476)(629,476){1}
wire w78;    //: /sn:0 {0}(-325,134)(-270,134)(-270,661)(323,661)(323,428)(519,428){1}
wire w10;    //: /sn:0 {0}(-325,34)(66,34)(66,93)(120,93){1}
wire w72;    //: /sn:0 {0}(519,524)(399,524)(399,801)(-178,801)(-178,634)(-325,634){1}
wire w13;    //: /sn:0 {0}(120,45)(106,45)(106,4)(-325,4){1}
wire w52;    //: /sn:0 {0}(-325,534)(-117,534)(-117,-59)(347,-59)(347,125)(519,125){1}
wire w33;    //: /sn:0 {0}(-325,104)(-238,104)(-238,451)(120,451){1}
wire w80;    //: /sn:0 {0}(614,524)(668,524){1}
wire w79;    //: /sn:0 {0}(-325,124)(-260,124)(-260,650)(314,650)(314,412)(519,412){1}
wire w50;    //: /sn:0 {0}(519,157)(324,157)(324,-33)(-90,-33)(-90,554)(-325,554){1}
wire w9;    //: /sn:0 {0}(120,109)(-204,109)(-204,484)(-325,484){1}
wire w55;    //: /sn:0 {0}(-325,64)(-157,64)(-157,-97)(383,-97)(383,77)(519,77){1}
wire w39;    //: /sn:0 {0}(215,483)(230,483){1}
//: enddecls

  //: OUT g4 (F) @(1045,256) /sn:0 /w:[ 0 ]
  //: joint g8 (w1) @(4, 275) /w:[ 9 -1 10 12 ]
  //: IN g3 (S) @(-408,290) /sn:0 /w:[ 0 ]
  //: joint g13 (w46) @(39, 285) /w:[ 3 4 6 -1 ]
  //: IN g2 (M) @(-408,368) /sn:0 /w:[ 13 ]
  //: IN g1 (B) @(-408,559) /sn:0 /w:[ 1 ]
  H74181 g11 (._A0(w35), ._A1(w34), ._A2(w33), ._A3(w32), ._B0(w31), ._B1(w30), ._B2(w40), ._B3(w28), .Cn(w60), .M(M), .S0(w1), .S1(w46), .S2(w45), .S3(w0), ._F0(w43), ._F1(w96), ._F2(w97), ._F3(w98), .AEB(w39), .CnP4(w38), ._G(w37), ._P(w36));   //: @(121, 403) /sz:(93, 240) /sn:0 /p:[ Li0>1 Li1>1 Li2>1 Li3>1 Li4>1 Li5>0 Li6>0 Li7>0 Li8>0 Li9>3 Li10>13 Li11>11 Li12>13 Li13>13 Ro0<0 Ro1<0 Ro2<0 Ro3<1 Ro4<0 Ro5<0 Ro6<0 Ro7<0 ]
  //: joint g16 (w1) @(233, 275) /w:[ 2 -1 4 1 ]
  assign {w76, w77, w78, w79, w32, w33, w34, w35, w54, w55, w56, w57, w10, w11, w12, w13} = A; //: CONCAT A_C  @(-330,79) /sn:0 /R:2 /w:[ 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 1 1 ] /dr:0 /tp:1 /drp:0
  H74181 g10 (._A0(w57), ._A1(w56), ._A2(w55), ._A3(w54), ._B0(w53), ._B1(w52), ._B2(w51), ._B3(w50), .Cn(w16), .M(M), .S0(w1), .S1(w46), .S2(w45), .S3(w0), ._F0(w65), ._F1(w64), ._F2(w93), ._F3(w62), .AEB(w61), .CnP4(w60), ._G(w59), ._P(w58));   //: @(520, 29) /sz:(93, 240) /sn:0 /p:[ Li0>1 Li1>1 Li2>1 Li3>1 Li4>0 Li5>1 Li6>1 Li7>0 Li8>1 Li9>9 Li10>3 Li11>0 Li12>3 Li13>3 Ro0<0 Ro1<0 Ro2<0 Ro3<0 Ro4<0 Ro5<1 Ro6<0 Ro7<0 ]
  //: joint g28 (w45) @(216, 295) /w:[ 2 -1 4 1 ]
  //: joint g19 (w0) @(207, 305) /w:[ 2 -1 4 1 ]
  //: joint g6 (M) @(18, 325) /w:[ 8 10 -1 7 ]
  H74181 g9 (._A0(w79), ._A1(w78), ._A2(w77), ._A3(w76), ._B0(w75), ._B1(w74), ._B2(w73), ._B3(w72), .Cn(w38), .M(M), .S0(w1), .S1(w46), .S2(w45), .S3(w0), ._F0(w99), ._F1(w100), ._F2(w101), ._F3(w102), .AEB(w83), .CnP4(CO), ._G(w81), ._P(w80));   //: @(520, 396) /sz:(93, 240) /sn:0 /p:[ Li0>1 Li1>1 Li2>0 Li3>0 Li4>0 Li5>0 Li6>0 Li7>0 Li8>1 Li9>0 Li10>0 Li11>13 Li12>0 Li13>0 Ro0<1 Ro1<0 Ro2<1 Ro3<0 Ro4<0 Ro5<1 Ro6<0 Ro7<0 ]
  //: joint g7 (w0) @(-27, 305) /w:[ 9 -1 10 12 ]
  //: joint g15 (w46) @(-6, 285) /w:[ 7 -1 8 10 ]
  //: IN g20 (CI) @(-408,218) /sn:0 /w:[ 1 ]
  //: joint g17 (M) @(18, 368) /w:[ -1 6 12 5 ]
  H74181 g29 (._A0(w13), ._A1(w12), ._A2(w11), ._A3(w10), ._B0(w9), ._B1(w8), ._B2(w7), ._B3(w6), .Cn(CI), .M(M), .S0(w1), .S1(w46), .S2(w45), .S3(w0), ._F0(w21), ._F1(w20), ._F2(w19), ._F3(w90), .AEB(w17), .CnP4(w16), ._G(w15), ._P(w14));   //: @(121, 29) /sz:(93, 240) /sn:0 /p:[ Li0>0 Li1>1 Li2>1 Li3>1 Li4>0 Li5>0 Li6>0 Li7>0 Li8>0 Li9>11 Li10>7 Li11>5 Li12>7 Li13>7 Ro0<0 Ro1<0 Ro2<0 Ro3<0 Ro4<0 Ro5<0 Ro6<0 Ro7<0 ]
  //: OUT g5 (CO) @(1022,491) /sn:0 /w:[ 0 ]
  assign {w0, w45, w46, w1} = S; //: CONCAT g14  @(-330,290) /sn:0 /R:2 /w:[ 11 11 9 11 1 ] /dr:0 /tp:1 /drp:0
  //: joint g24 (M) @(19, 563) /w:[ 2 4 -1 1 ]
  //: joint g21 (w46) @(225, 285) /w:[ 1 -1 2 12 ]
  assign F = {w102, w101, w100, w99, w98, w97, w96, w43, w62, w93, w64, w65, w90, w19, w20, w21}; //: CONCAT g23  @(985,256) /sn:0 /w:[ 1 1 0 1 0 0 1 1 1 1 1 1 1 1 1 1 1 ] /dr:1 /tp:1 /drp:1
  //: IN g0 (A) @(-408,79) /sn:0 /w:[ 0 ]
  //: joint g22 (w45) @(48, 295) /w:[ 5 6 8 -1 ]
  assign {w72, w73, w74, w75, w28, w40, w30, w31, w50, w51, w52, w53, w6, w7, w8, w9} = B; //: CONCAT B_C  @(-330,559) /sn:0 /R:2 /w:[ 1 1 1 1 1 1 1 0 1 0 0 1 1 1 1 1 0 ] /dr:0 /tp:0 /drp:0
  //: joint g12 (w45) @(-17, 295) /w:[ 9 -1 10 12 ]
  //: joint g18 (w0) @(57, 305) /w:[ 5 6 8 -1 ]
  //: joint g30 (w1) @(29, 275) /w:[ 5 6 8 -1 ]

endmodule
//: /netlistEnd

//: /netlistBegin ALU16_74181_74182
module ALU16_74181_74182(CI, F, OP, B, M, CO, A);
//: interface  /sz:(196, 96) /bd:[ Li0>A[15:0](16/96) Li1>B[15:0](32/96) Li2>CI(48/96) Li3>M(64/96) Li4>OP[3:0](80/96) Ro0<CO(16/96) Ro1<F[15:0](32/96) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input M;    //: /sn:0 {0}(630,91)(536,91)(536,183)(303,183){1}
//: {2}(301,181)(301,87)(351,87){3}
//: {4}(299,183)(173,183)(173,183)(49,183){5}
input [15:0] B;    //: /sn:0 {0}(#:50:98,355)(72,355)(72,355)(#:49,355){1}
output [15:0] F;    //: /sn:0 {0}(#:812,247)(827,247){1}
input [15:0] A;    //: /sn:0 {0}(#:49,18)(74,18)(74,18)(#:98,18){1}
output CO;    //: /sn:0 {0}(812,360)(827,360){1}
input [3:0] OP;    //: /sn:0 {0}(#:54,495)(#:95,495){1}
input CI;    //: /sn:0 {0}(351,71)(315,71)(315,373){1}
//: {2}(313,375)(164,375){3}
//: {4}(315,377)(315,571)(598,571){5}
wire w6;    //: /sn:0 {0}(598,475)(583,475){1}
wire w32;    //: /sn:0 {0}(446,-25)(461,-25){1}
wire w7;    //: /sn:0 {0}(725,43)(827,43)(827,215)(580,215)(580,459)(598,459){1}
wire w45;    //: /sn:0 {0}(104,-17)(208,-17)(208,-119)(612,-119)(612,-53)(630,-53){1}
wire w73;    //: /sn:0 {0}(104,400)(119,400){1}
wire w46;    //: /sn:0 {0}(725,59)(815,59)(815,204)(577,204)(577,523)(598,523){1}
wire w61;    //: /sn:0 {0}(104,23)(119,23){1}
wire w14;    //: /sn:0 {0}(351,135)(205,135)(205,500)(101,500){1}
wire w4;    //: /sn:0 {0}(598,507)(463,507)(463,55)(446,55){1}
wire w15;    //: /sn:0 {0}(630,123)(559,123)(559,420){1}
//: {2}(557,422)(197,422){3}
//: {4}(195,420)(195,119)(351,119){5}
//: {6}(195,424)(195,490)(101,490){7}
//: {8}(559,424)(559,431){9}
wire w19;    //: /sn:0 {0}(351,55)(291,55)(291,310)(104,310){1}
wire w38;    //: /sn:0 {0}(630,59)(525,59)(525,350)(104,350){1}
wire w51;    //: /sn:0 {0}(725,-21)(740,-21){1}
wire w69;    //: /sn:0 {0}(104,360)(119,360){1}
wire w3;    //: /sn:0 {0}(351,103)(183,103)(183,403){1}
//: {2}(185,405)(549,405)(549,107)(630,107){3}
//: {4}(183,407)(183,480)(101,480){5}
wire w0;    //: /sn:0 {0}(351,151)(218,151)(218,510)(101,510){1}
wire w37;    //: /sn:0 {0}(630,75)(615,75){1}
wire w64;    //: /sn:0 {0}(104,53)(119,53){1}
wire w66;    //: /sn:0 {0}(104,73)(119,73){1}
wire w34;    //: /sn:0 {0}(446,-57)(461,-57){1}
wire w63;    //: /sn:0 {0}(104,43)(119,43){1}
wire w21;    //: /sn:0 {0}(104,290)(268,290)(268,23)(351,23){1}
wire w43;    //: /sn:0 {0}(630,-21)(586,-21)(586,-92)(231,-92)(231,3)(104,3){1}
wire w75;    //: /sn:0 {0}(104,420)(119,420){1}
wire w76;    //: /sn:0 {0}(104,430)(119,430){1}
wire w67;    //: /sn:0 {0}(104,83)(119,83){1}
wire w31;    //: /sn:0 {0}(446,-9)(461,-9){1}
wire w58;    //: /sn:0 {0}(630,43)(512,43)(512,340)(104,340){1}
wire w20;    //: /sn:0 {0}(351,39)(280,39)(280,300)(104,300){1}
wire w23;    //: /sn:0 {0}(104,-27)(271,-27)(271,-9)(351,-9){1}
wire w24;    //: /sn:0 {0}(104,-37)(280,-37)(280,-25)(351,-25){1}
wire w41;    //: /sn:0 {0}(630,11)(487,11)(487,320)(104,320){1}
wire w1;    //: /sn:0 {0}(598,555)(583,555){1}
wire w25;    //: /sn:0 {0}(104,-47)(292,-47)(292,-41)(351,-41){1}
wire w65;    //: /sn:0 {0}(104,63)(119,63){1}
wire w74;    //: /sn:0 {0}(104,410)(119,410){1}
wire w8;    //: /sn:0 {0}(598,443)(474,443)(474,39)(446,39){1}
wire w18;    //: /sn:0 {0}(630,155)(615,155){1}
wire w40;    //: /sn:0 {0}(630,27)(499,27)(499,330)(104,330){1}
wire w30;    //: /sn:0 {0}(446,7)(461,7){1}
wire w68;    //: /sn:0 {0}(104,93)(119,93){1}
wire w71;    //: /sn:0 {0}(104,380)(119,380){1}
wire w22;    //: /sn:0 {0}(351,7)(258,7)(258,280)(104,280){1}
wire w53;    //: /sn:0 {0}(725,-53)(740,-53){1}
wire w62;    //: /sn:0 {0}(104,33)(119,33){1}
wire w2;    //: /sn:0 {0}(598,539)(583,539){1}
wire w11;    //: /sn:0 {0}(705,475)(720,475){1}
wire w12;    //: /sn:0 {0}(705,459)(720,459){1}
wire w44;    //: /sn:0 {0}(630,-37)(600,-37)(600,-106)(219,-106)(219,-7)(104,-7){1}
wire w49;    //: /sn:0 {0}(725,11)(740,11){1}
wire w70;    //: /sn:0 {0}(104,370)(119,370){1}
wire w10;    //: /sn:0 {0}(705,491)(720,491){1}
wire w13;    //: /sn:0 {0}(705,443)(720,443){1}
wire w27;    //: /sn:0 {0}(630,139)(615,139){1}
wire w72;    //: /sn:0 {0}(104,390)(119,390){1}
wire w5;    //: /sn:0 {0}(598,491)(583,491){1}
wire w33;    //: /sn:0 {0}(446,-41)(461,-41){1}
wire w48;    //: /sn:0 {0}(725,27)(740,27){1}
wire w52;    //: /sn:0 {0}(725,-37)(740,-37){1}
wire w29;    //: /sn:0 {0}(446,23)(461,23){1}
wire w9;    //: /sn:0 {0}(705,507)(720,507){1}
wire w42;    //: /sn:0 {0}(630,-5)(573,-5)(573,-78)(244,-78)(244,13)(104,13){1}
wire w50;    //: /sn:0 {0}(725,-5)(740,-5){1}
wire w26;    //: /sn:0 {0}(104,-57)(351,-57){1}
//: enddecls

  //: IN g4 (CI) @(162,375) /sn:0 /w:[ 3 ]
  H74181 g8 (._A0(w26), ._A1(w25), ._A2(w24), ._A3(w23), ._B0(w22), ._B1(w21), ._B2(w20), ._B3(w19), .Cn(CI), .M(M), .S0(w3), .S1(w15), .S2(w14), .S3(w0), ._F0(w34), ._F1(w33), ._F2(w32), ._F3(w31), .AEB(w30), .CnP4(w29), ._G(w8), ._P(w4));   //: @(352, -73) /sz:(93, 240) /sn:0 /p:[ Li0>1 Li1>1 Li2>1 Li3>1 Li4>0 Li5>1 Li6>0 Li7>0 Li8>0 Li9>3 Li10>0 Li11>5 Li12>0 Li13>0 Ro0<0 Ro1<0 Ro2<0 Ro3<0 Ro4<0 Ro5<0 Ro6<1 Ro7<1 ]
  //: OUT g3 (F) @(824,247) /sn:0 /w:[ 1 ]
  assign {w76, w75, w74, w73, w72, w71, w70, w69, w38, w58, w40, w41, w19, w20, w21, w22} = B; //: CONCAT g13  @(99,355) /sn:0 /R:2 /w:[ 0 0 0 0 0 0 0 0 1 1 1 1 1 1 0 1 0 ] /dr:0 /tp:1 /drp:0
  //: IN g2 (OP) @(52,495) /sn:0 /w:[ 0 ]
  //: IN g1 (B) @(47,355) /sn:0 /w:[ 1 ]
  //: joint g16 (w3) @(183, 405) /w:[ 2 1 -1 4 ]
  assign {w68, w67, w66, w65, w64, w63, w62, w61, w42, w43, w44, w45, w23, w24, w25, w26} = A; //: CONCAT g11  @(99,18) /sn:0 /R:2 /w:[ 0 0 0 0 0 0 0 0 1 1 1 0 0 0 0 0 1 ] /dr:0 /tp:1 /drp:0
  H74181 g10 (._A0(w45), ._A1(w44), ._A2(w43), ._A3(w42), ._B0(w41), ._B1(w40), ._B2(w58), ._B3(w38), .Cn(w37), .M(M), .S0(w3), .S1(w15), .S2(w27), .S3(w18), ._F0(w53), ._F1(w52), ._F2(w51), ._F3(w50), .AEB(w49), .CnP4(w48), ._G(w7), ._P(w46));   //: @(631, -69) /sz:(93, 240) /sn:0 /p:[ Li0>1 Li1>0 Li2>0 Li3>0 Li4>0 Li5>0 Li6>0 Li7>0 Li8>0 Li9>0 Li10>3 Li11>0 Li12>0 Li13>0 Ro0<0 Ro1<0 Ro2<0 Ro3<0 Ro4<0 Ro5<0 Ro6<0 Ro7<0 ]
  //: IN g6 (M) @(47,183) /sn:0 /w:[ 5 ]
  H74182 g7 (._G0(w8), ._G1(w7), ._G2(w6), ._G3(w5), ._P0(w4), ._P1(w46), ._P2(w2), ._P3(w1), .Cn(CI), .CnPx(w13), .CnPy(w12), .CnPz(w11), ._G(w10), ._P(w9));   //: @(599, 427) /sz:(105, 160) /sn:0 /p:[ Li0>0 Li1>1 Li2>0 Li3>0 Li4>0 Li5>1 Li6>0 Li7>0 Li8>5 Ro0<0 Ro1<0 Ro2<0 Ro3<0 Ro4<0 ]
  //: joint g9 (CI) @(315, 375) /w:[ -1 1 2 4 ]
  //: joint g15 (w15) @(559, 422) /w:[ -1 1 2 8 ]
  //: joint g17 (w15) @(195, 422) /w:[ 3 4 -1 6 ]
  assign {w0, w14, w15, w3} = OP; //: CONCAT g14  @(96,495) /sn:0 /R:2 /w:[ 1 1 7 5 1 ] /dr:0 /tp:0 /drp:0
  //: OUT g5 (CO) @(824,360) /sn:0 /w:[ 1 ]
  //: IN g0 (A) @(47,18) /sn:0 /w:[ 0 ]
  //: joint g12 (M) @(301, 183) /w:[ 1 2 4 -1 ]

endmodule
//: /netlistEnd


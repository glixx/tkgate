//: version "2.0-b10"
//: property encoding = "utf-8"
//: property locale = "ru"
//: property prefix = "_GG"
//: property title = "Микросхемы стандартной логики"
//: property timingViolationMode = 2
//: property initTime = "0 ns"
//: require "74xx"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg [15:0] A_NET;    //: {0}(#:79,174)(144,174)(144,174)(213,174){1}
//: {2}(1:217,174)(271,174){3}
//: {4}(#:215,176)(215,352)(268,352){5}
reg [3:0] OP_NET;    //: {0}(#:78,417)(114,417){1}
//: {2}(-18:118,417)(193,417)(193,416)(268,416){3}
//: {4}(116,415)(116,238)(271,238){5}
reg w0;    //: /sn:0 {0}(56,380)(149,380){1}
//: {2}(151,378)(151,222)(271,222){3}
//: {4}(151,382)(151,400)(268,400){5}
reg w3;    //: /sn:0 {0}(58,323)(163,323){1}
//: {2}(165,321)(165,206)(271,206){3}
//: {4}(165,325)(165,384)(268,384){5}
reg [15:0] B_NET;    //: {0}(#:79,228)(102,228)(64:102,190)(178,190){1}
//: {2}(182,190)(271,190){3}
//: {4}(#:180,192)(180,368)(268,368){5}
wire [15:0] pulse;    //: /sn:0 {0}(#:513,190)(415,190){1}
wire [15:0] propagation;    //: /sn:0 {0}(#:513,369)(490,369)(490,368)(466,368){1}
wire w11;    //: /sn:0 {0}(479,325)(479,352)(466,352){1}
wire w5;    //: /sn:0 {0}(415,174)(479,174)(479,148){1}
//: enddecls

  //: SWITCH M (w0) @(39,380) /w:[ 0 ] /st:0 /dn:1
  //: joint g4 (A_NET) @(215, 174) /w:[ 2 -1 1 4 ]
  //: joint g8 (w0) @(151, 380) /w:[ -1 2 1 4 ]
  ALU16_74181_74182 g3 (.A(A_NET), .B(B_NET), .CI(w3), .M(w0), .OP(OP_NET), .CO(w11), .F(propagation));   //: @(269, 336) /sz:(196, 96) /sn:0 /p:[ Li0>5 Li1>5 Li2>5 Li3>5 Li4>3 Ro0<1 Ro1<1 ]
  //: comment g2 @(74,9) /sn:0
  //: /line:"     Логические (M=1)"
  //: /line:"00 - НЕ <b>A</b>"
  //: /line:"01 - <b>A</b> НЕ-ИЛИ <b>B</b>"
  //: /line:"02 - НЕ <b>A</b> И <b>B</b>"
  //: /line:"05 - НЕ <b>B</b>"
  //: /line:"06 - <b>A</b> ИСКЛ. ИЛИ <b>B</b>"
  //: /line:"09 - <b>A</b> НЕ-ИСКЛ. ИЛИ <b>B</b>"
  //: /line:"0B - <b>A</b> И <b>B</b>"
  //: /line:"0E - <b>A</b> ИЛИ <b>B</b>"
  //: /end
  //: LED g1 (w5) @(479,141) /sn:0 /w:[ 1 ] /type:0
  //: DIP B_DIP (B_NET) @(41,228) /R:1 /w:[ 0 ] /st:2 /dn:1
  //: DIP OP_DIP (OP_NET) @(40,417) /R:1 /w:[ 0 ] /st:1 /dn:1
  //: LED g11 (propagation) @(520,369) /sn:0 /R:3 /w:[ 0 ] /type:2
  //: LED g10 (w11) @(479,318) /sn:0 /w:[ 0 ] /type:0
  //: LED g6 (pulse) @(520,190) /sn:0 /R:3 /w:[ 0 ] /type:2
  //: joint g7 (w3) @(165, 323) /w:[ -1 2 1 4 ]
  //: joint g9 (OP_NET) @(116, 417) /w:[ 2 4 1 -1 ]
  //: SWITCH CI (w3) @(41,323) /w:[ 0 ] /st:1 /dn:1
  //: joint g5 (B_NET) @(180, 190) /w:[ 2 -1 1 4 ]
  ALU16_74181 g0 (.A(A_NET), .B(B_NET), .CI(w3), .M(w0), .S(OP_NET), .CO(w5), .F(pulse));   //: @(272, 158) /sz:(142, 96) /sn:0 /p:[ Li0>3 Li1>3 Li2>3 Li3>3 Li4>5 Ro0<0 Ro1<1 ]
  //: DIP A_DIP (A_NET) @(41,174) /R:1 /w:[ 0 ] /st:2 /dn:1
  //: comment g12 @(210,9) /sn:0
  //: /line:"  Арифметические (M=0)"
  //: /line:"<b>A</b>"
  //: /line:"<b>A</b> ИЛИ <b>B</b>"
  //: /line:"<b>A</b> ИЛИ НЕ <b>B</b>"
  //: /line:"(<b>A</b> ИЛИ <b>B</b>)+(<b>A</b> И НЕ <b>B</b>)"
  //: /line:"<b>A</b> - <b>B</b> - 1"
  //: /line:"<b>A</b> + <b>B</b>"
  //: /line:"<b>A</b> И <b>B</b> - 1"
  //: /line:"<b>A</b> ИЛИ <b>B</b>"
  //: /end

endmodule
//: /netlistEnd

//: /netlistBegin ALU16_74181
module ALU16_74181(F, S, M, B, CI, CO, A);
//: interface  /sz:(142, 96) /bd:[ Li0>A[15:0](16/96) Li1>B[15:0](32/96) Li2>CI(48/96) Li3>M(64/96) Li4>S[3:0](80/96) Ro0<CO(16/96) Ro1<F[15:0](32/96) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input M;    //: {0}(519,556)(353,556)(353,695)(19,695)(19,565){1}
//: {2}(21,563)(71,563)(71,563)(120,563){3}
//: {4}(19,561)(19,465)(18,465)(18,370){5}
//: {6}(18,366)(18,327){7}
//: {8}(20,325)(429,325)(429,189)(519,189){9}
//: {10}(18,323)(18,189)(120,189){11}
//: {12}(16,368)(-194,368)(-194,368)(99:-406,368){13}
input [15:0] B;    //: /sn:0 {0}(#:-331,559)(#:-406,559){1}
output [15:0] F;    //: /sn:0 {0}(1048,256)(#:986,256){1}
input [15:0] A;    //: {0}(#:80:-406,79)(-373,79)(-373,79)(#:58:-331,79){1}
output CO;    //: /sn:0 {0}(1025,491)(819,491)(819,492)(614,492){1}
input CI;    //: /sn:0 {0}(120,173)(-347,173)(-347,218)(-406,218){1}
input [3:0] S;    //: {0}(#:70:-406,290)(-367,290)(-367,290)(#:-331,290){1}
wire w32;    //: /sn:0 {0}(-325,114)(-249,114)(-249,467)(120,467){1}
wire w6;    //: /sn:0 {0}(120,157)(-171,157)(-171,514)(-325,514){1}
wire w73;    //: /sn:0 {0}(519,508)(386,508)(386,789)(-169,789)(-169,624)(-325,624){1}
wire w45;    //: /sn:0 {0}(519,604)(471,604)(471,355)(216,355)(216,297){1}
//: {2}(218,295)(466,295)(466,237)(519,237){3}
//: {4}(214,295)(50,295){5}
//: {6}(48,293)(48,237)(120,237){7}
//: {8}(46,295)(-15,295){9}
//: {10}(-19,295)(-325,295){11}
//: {12}(-17,297)(-17,611)(120,611){13}
wire w93;    //: /sn:0 {0}(614,77)(906,77)(906,241)(980,241){1}
wire w96;    //: /sn:0 {0}(215,435)(288,435)(288,736)(863,736)(863,271)(980,271){1}
wire w7;    //: /sn:0 {0}(120,141)(-182,141)(-182,504)(-325,504){1}
wire w46;    //: /sn:0 {0}(519,221)(453,221)(453,285)(227,285){1}
//: {2}(223,285)(41,285){3}
//: {4}(39,283)(39,221)(120,221){5}
//: {6}(37,285)(-4,285){7}
//: {8}(-8,285)(-325,285){9}
//: {10}(-6,287)(-6,595)(120,595){11}
//: {12}(225,287)(225,346)(481,346)(481,588)(519,588){13}
wire w99;    //: /sn:0 {0}(980,301)(893,301)(893,412)(614,412){1}
wire w61;    //: /sn:0 {0}(614,109)(629,109){1}
wire w60;    //: /sn:0 {0}(120,547)(35,547)(35,706)(841,706)(841,125)(614,125){1}
wire w56;    //: /sn:0 {0}(519,61)(490,61)(490,63)(475,63){1}
wire w16;    //: /sn:0 {0}(215,125)(310,125)(310,173)(519,173){1}
wire w14;    //: /sn:0 {0}(215,157)(230,157){1}
wire w81;    //: /sn:0 {0}(614,508)(629,508){1}
wire w19;    //: /sn:0 {0}(215,77)(297,77)(297,6)(945,6)(945,201)(980,201){1}
wire w15;    //: /sn:0 {0}(215,141)(230,141){1}
wire w38;    //: /sn:0 {0}(215,499)(251,499)(251,540)(519,540){1}
wire w51;    //: /sn:0 {0}(-325,544)(-104,544)(-104,-46)(336,-46)(336,141)(519,141){1}
wire w0;    //: /sn:0 {0}(519,620)(460,620)(460,363)(207,363)(207,307){1}
//: {2}(209,305)(478,305)(478,253)(519,253){3}
//: {4}(205,305)(59,305){5}
//: {6}(57,303)(57,253)(120,253){7}
//: {8}(55,305)(-25,305){9}
//: {10}(-29,305)(-325,305){11}
//: {12}(-27,307)(-27,627)(120,627){13}
wire w97;    //: /sn:0 {0}(215,451)(277,451)(277,747)(875,747)(875,281)(980,281){1}
wire w3;    //: /sn:0 {0}(-273,54)(-325,54){1}
wire w64;    //: /sn:0 {0}(614,61)(917,61)(917,231)(980,231){1}
wire w37;    //: /sn:0 {0}(215,515)(230,515){1}
wire w34;    //: /sn:0 {0}(-325,94)(-227,94)(-227,435)(120,435){1}
wire w76;    //: /sn:0 {0}(519,460)(343,460)(343,683)(-288,683)(-288,154)(-325,154){1}
wire w75;    //: /sn:0 {0}(519,476)(363,476)(363,765)(-148,765)(-148,604)(-325,604){1}
wire w102;    //: /sn:0 {0}(614,460)(922,460)(922,331)(980,331){1}
wire w43;    //: /sn:0 {0}(215,419)(299,419)(299,726)(851,726)(851,261)(980,261){1}
wire w21;    //: /sn:0 {0}(215,45)(273,45)(273,-19)(966,-19)(966,181)(980,181){1}
wire w54;    //: /sn:0 {0}(519,93)(490,93)(490,83)(475,83){1}
wire w100;    //: /sn:0 {0}(614,428)(902,428)(902,311)(980,311){1}
wire w58;    //: /sn:0 {0}(614,157)(629,157){1}
wire w31;    //: /sn:0 {0}(-325,564)(-77,564)(-77,483)(120,483){1}
wire w90;    //: /sn:0 {0}(215,93)(308,93)(308,21)(934,21)(934,211)(980,211){1}
wire w28;    //: /sn:0 {0}(120,531)(-39,531)(-39,594)(-325,594){1}
wire w36;    //: /sn:0 {0}(215,531)(230,531){1}
wire w20;    //: /sn:0 {0}(215,61)(285,61)(285,-6)(956,-6)(956,191)(980,191){1}
wire w1;    //: /sn:0 {0}(519,572)(490,572)(490,336)(233,336)(233,277){1}
//: {2}(235,275)(441,275)(441,205)(519,205){3}
//: {4}(231,275)(31,275){5}
//: {6}(29,273)(29,205)(120,205){7}
//: {8}(27,275)(6,275){9}
//: {10}(2,275)(-325,275){11}
//: {12}(4,277)(4,579)(120,579){13}
wire w74;    //: /sn:0 {0}(519,492)(374,492)(374,776)(-159,776)(-159,614)(-325,614){1}
wire w65;    //: /sn:0 {0}(614,45)(926,45)(926,221)(980,221){1}
wire w98;    //: /sn:0 {0}(980,291)(887,291)(887,756)(264,756)(264,467)(215,467){1}
wire w40;    //: /sn:0 {0}(120,515)(-50,515)(-50,584)(-325,584){1}
wire w35;    //: /sn:0 {0}(-325,84)(-215,84)(-215,419)(120,419){1}
wire w8;    //: /sn:0 {0}(120,125)(-195,125)(-195,494)(-325,494){1}
wire w18;    //: /sn:0 {0}(-273,74)(-325,74){1}
wire w101;    //: /sn:0 {0}(980,321)(912,321)(912,444)(614,444){1}
wire w30;    //: /sn:0 {0}(120,499)(-64,499)(-64,574)(-325,574){1}
wire w17;    //: /sn:0 {0}(215,109)(230,109){1}
wire [3:0] w22;    //: /sn:0 {0}(#:469,68)(431,68)(431,-90)(-226,-90)(-226,59)(#:-267,59){1}
wire w53;    //: /sn:0 {0}(519,109)(358,109)(358,-72)(-130,-72)(-130,524)(-325,524){1}
wire w59;    //: /sn:0 {0}(614,141)(629,141){1}
wire w62;    //: /sn:0 {0}(614,93)(897,93)(897,251)(980,251){1}
wire w57;    //: /sn:0 {0}(519,45)(490,45)(490,53)(475,53){1}
wire w12;    //: /sn:0 {0}(-325,14)(94,14)(94,61)(120,61){1}
wire w11;    //: /sn:0 {0}(-325,24)(80,24)(80,77)(120,77){1}
wire w2;    //: /sn:0 {0}(-273,44)(-325,44){1}
wire w77;    //: /sn:0 {0}(519,444)(333,444)(333,672)(-279,672)(-279,144)(-325,144){1}
wire w83;    //: /sn:0 {0}(614,476)(629,476){1}
wire w78;    //: /sn:0 {0}(-325,134)(-270,134)(-270,661)(323,661)(323,428)(519,428){1}
wire w10;    //: /sn:0 {0}(-325,34)(66,34)(66,93)(120,93){1}
wire w72;    //: /sn:0 {0}(519,524)(399,524)(399,801)(-178,801)(-178,634)(-325,634){1}
wire w13;    //: /sn:0 {0}(120,45)(106,45)(106,4)(-325,4){1}
wire w52;    //: /sn:0 {0}(-325,534)(-117,534)(-117,-59)(347,-59)(347,125)(519,125){1}
wire w33;    //: /sn:0 {0}(-325,104)(-238,104)(-238,451)(120,451){1}
wire w5;    //: /sn:0 {0}(-273,64)(-325,64){1}
wire w80;    //: /sn:0 {0}(614,524)(668,524){1}
wire w79;    //: /sn:0 {0}(-325,124)(-260,124)(-260,650)(314,650)(314,412)(519,412){1}
wire w50;    //: /sn:0 {0}(519,157)(324,157)(324,-33)(-90,-33)(-90,554)(-325,554){1}
wire w9;    //: /sn:0 {0}(120,109)(-204,109)(-204,484)(-325,484){1}
wire w55;    //: /sn:0 {0}(519,77)(490,77)(490,73)(475,73){1}
wire w39;    //: /sn:0 {0}(215,483)(230,483){1}
//: enddecls

  //: OUT g4 (F) @(1045,256) /sn:0 /w:[ 0 ]
  //: joint g8 (w1) @(4, 275) /w:[ 9 -1 10 12 ]
  //: IN g3 (S) @(-408,290) /sn:0 /w:[ 0 ]
  //: joint g13 (w46) @(39, 285) /w:[ 3 4 6 -1 ]
  //: IN g2 (M) @(-408,368) /sn:0 /w:[ 13 ]
  //: IN g1 (B) @(-408,559) /sn:0 /w:[ 1 ]
  H74181 g11 (._A0(w35), ._A1(w34), ._A2(w33), ._A3(w32), ._B0(w31), ._B1(w30), ._B2(w40), ._B3(w28), .Cn(w60), .M(M), .S0(w1), .S1(w46), .S2(w45), .S3(w0), ._F0(w43), ._F1(w96), ._F2(w97), ._F3(w98), .AEB(w39), .CnP4(w38), ._G(w37), ._P(w36));   //: @(121, 403) /sz:(93, 240) /sn:0 /p:[ Li0>1 Li1>1 Li2>1 Li3>1 Li4>1 Li5>0 Li6>0 Li7>0 Li8>0 Li9>3 Li10>13 Li11>11 Li12>13 Li13>13 Ro0<0 Ro1<0 Ro2<0 Ro3<1 Ro4<0 Ro5<0 Ro6<0 Ro7<0 ]
  //: joint g16 (w1) @(233, 275) /w:[ 2 -1 4 1 ]
  assign {w76, w77, w78, w79, w32, w33, w34, w35, w18, w5, w3, w2, w10, w11, w12, w13} = A; //: CONCAT A_C  @(-330,79) /sn:0 /R:2 /w:[ 1 1 0 0 0 0 0 0 1 1 1 1 0 0 0 1 1 ] /dr:0 /tp:1 /drp:0
  H74181 g10 (._A0(w57), ._A1(w56), ._A2(w55), ._A3(w54), ._B0(w53), ._B1(w52), ._B2(w51), ._B3(w50), .Cn(w16), .M(M), .S0(w1), .S1(w46), .S2(w45), .S3(w0), ._F0(w65), ._F1(w64), ._F2(w93), ._F3(w62), .AEB(w61), .CnP4(w60), ._G(w59), ._P(w58));   //: @(520, 29) /sz:(93, 240) /sn:0 /p:[ Li0>0 Li1>0 Li2>0 Li3>0 Li4>0 Li5>1 Li6>1 Li7>0 Li8>1 Li9>9 Li10>3 Li11>0 Li12>3 Li13>3 Ro0<0 Ro1<0 Ro2<0 Ro3<0 Ro4<0 Ro5<1 Ro6<0 Ro7<0 ]
  //: joint g28 (w45) @(216, 295) /w:[ 2 -1 4 1 ]
  //: joint g19 (w0) @(207, 305) /w:[ 2 -1 4 1 ]
  //: joint g6 (M) @(18, 325) /w:[ 8 10 -1 7 ]
  H74181 g9 (._A0(w79), ._A1(w78), ._A2(w77), ._A3(w76), ._B0(w75), ._B1(w74), ._B2(w73), ._B3(w72), .Cn(w38), .M(M), .S0(w1), .S1(w46), .S2(w45), .S3(w0), ._F0(w99), ._F1(w100), ._F2(w101), ._F3(w102), .AEB(w83), .CnP4(CO), ._G(w81), ._P(w80));   //: @(520, 396) /sz:(93, 240) /sn:0 /p:[ Li0>1 Li1>1 Li2>0 Li3>0 Li4>0 Li5>0 Li6>0 Li7>0 Li8>1 Li9>0 Li10>0 Li11>13 Li12>0 Li13>0 Ro0<1 Ro1<0 Ro2<1 Ro3<0 Ro4<0 Ro5<1 Ro6<0 Ro7<0 ]
  //: joint g7 (w0) @(-27, 305) /w:[ 9 -1 10 12 ]
  //: joint g15 (w46) @(-6, 285) /w:[ 7 -1 8 10 ]
  //: IN g20 (CI) @(-408,218) /sn:0 /w:[ 1 ]
  //: joint g17 (M) @(18, 368) /w:[ -1 6 12 5 ]
  H74181 g29 (._A0(w13), ._A1(w12), ._A2(w11), ._A3(w10), ._B0(w9), ._B1(w8), ._B2(w7), ._B3(w6), .Cn(CI), .M(M), .S0(w1), .S1(w46), .S2(w45), .S3(w0), ._F0(w21), ._F1(w20), ._F2(w19), ._F3(w90), .AEB(w17), .CnP4(w16), ._G(w15), ._P(w14));   //: @(121, 29) /sz:(93, 240) /sn:0 /p:[ Li0>0 Li1>1 Li2>1 Li3>1 Li4>0 Li5>0 Li6>0 Li7>0 Li8>0 Li9>11 Li10>7 Li11>5 Li12>7 Li13>7 Ro0<0 Ro1<0 Ro2<0 Ro3<0 Ro4<0 Ro5<0 Ro6<0 Ro7<0 ]
  assign w22 = {w18, w5, w3, w2}; //: CONCAT g25  @(-268,59) /sn:0 /w:[ 1 0 0 0 0 ] /dr:1 /tp:1 /drp:1
  //: OUT g5 (CO) @(1022,491) /sn:0 /w:[ 0 ]
  assign {w0, w45, w46, w1} = S; //: CONCAT g14  @(-330,290) /sn:0 /R:2 /w:[ 11 11 9 11 1 ] /dr:0 /tp:1 /drp:0
  //: joint g24 (M) @(19, 563) /w:[ 2 4 -1 1 ]
  //: joint g21 (w46) @(225, 285) /w:[ 1 -1 2 12 ]
  assign F = {w102, w101, w100, w99, w98, w97, w96, w43, w62, w93, w64, w65, w90, w19, w20, w21}; //: CONCAT g23  @(985,256) /sn:0 /w:[ 1 1 0 1 0 0 1 1 1 1 1 1 1 1 1 1 1 ] /dr:1 /tp:1 /drp:1
  //: IN g0 (A) @(-408,79) /sn:0 /w:[ 0 ]
  //: joint g22 (w45) @(48, 295) /w:[ 5 6 8 -1 ]
  assign {w54, w55, w56, w57} = w22; //: CONCAT g26  @(470,68) /sn:0 /R:2 /w:[ 1 1 1 1 0 ] /dr:0 /tp:1 /drp:0
  assign {w72, w73, w74, w75, w28, w40, w30, w31, w50, w51, w52, w53, w6, w7, w8, w9} = B; //: CONCAT B_C  @(-330,559) /sn:0 /R:2 /w:[ 1 1 1 1 1 1 1 0 1 0 0 1 1 1 1 1 0 ] /dr:0 /tp:0 /drp:0
  //: joint g12 (w45) @(-17, 295) /w:[ 9 -1 10 12 ]
  //: joint g18 (w0) @(57, 305) /w:[ 5 6 8 -1 ]
  //: joint g30 (w1) @(29, 275) /w:[ 5 6 8 -1 ]

endmodule
//: /netlistEnd

//: /netlistBegin ALU16_74181_74182
module ALU16_74181_74182(CI, F, OP, B, M, CO, A);
//: interface  /sz:(196, 96) /bd:[ Li0>A[15:0](16/96) Li1>B[15:0](32/96) Li2>CI(48/96) Li3>M(64/96) Li4>OP[3:0](80/96) Ro0<CO(16/96) Ro1<F[15:0](32/96) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input M;    //: /sn:0 {0}(689,368)(571,368)(571,185){1}
//: {2}(571,181)(571,90)(689,90){3}
//: {4}(569,183)(314,183){5}
//: {6}(312,181)(312,87)(351,87){7}
//: {8}(310,183)(14,183){9}
//: {10}(312,185)(312,380)(347,380){11}
input [15:0] A;    //: /sn:0 {0}(#:14,18)(39,18)(39,18)(#:63,18){1}
output CO;    //: /sn:0 {0}(994,307)(799,307)(799,304)(784,304){1}
input [15:0] B;    //: /sn:0 {0}(#:50:105,553)(79,553)(79,553)(#:56,553){1}
output [15:0] F;    //: /sn:0 {0}(#:1017,62)(1053,62){1}
input [3:0] OP;    //: /sn:0 {0}(#:628,411)(595,411)(595,211){1}
//: {2}(595,207)(595,130)(#:628,130){3}
//: {4}(593,209)(220,209){5}
//: {6}(218,207)(218,127)(#:242,127){7}
//: {8}(216,209)(#:19,209){9}
//: {10}(218,211)(218,421)(#:247,421){11}
input CI;    //: /sn:0 {0}(351,71)(325,71)(325,655){1}
//: {2}(323,657)(135,657)(135,658)(58,658){3}
//: {4}(325,659)(325,771)(727,771){5}
wire w32;    //: /sn:0 {0}(488,-28)(457,-28)(457,-25)(446,-25){1}
wire w45;    //: /sn:0 {0}(689,-54)(649,-54)(649,-42)(634,-42){1}
wire w73;    //: /sn:0 {0}(153,599)(118,599)(118,598)(111,598){1}
wire w96;    //: /sn:0 {0}(634,308)(662,308)(662,304)(689,304){1}
wire [3:0] w16;    //: /sn:0 {0}(#:628,313)(550,313)(550,614)(#:159,614){1}
wire [3:0] w14;    //: /sn:0 {0}(#:125,78)(150,78)(150,199)(607,199)(607,252)(#:628,252){1}
wire w56;    //: /sn:0 {0}(916,67)(1011,67){1}
wire w4;    //: /sn:0 {0}(727,707)(507,707)(507,55)(446,55){1}
wire w19;    //: /sn:0 {0}(351,55)(298,55)(298,508)(111,508){1}
wire w89;    //: /sn:0 {0}(481,275)(472,275)(472,284)(442,284){1}
wire w81;    //: /sn:0 {0}(634,237)(643,237)(643,224)(689,224){1}
wire w38;    //: /sn:0 {0}(153,547)(113,547)(113,548)(111,548){1}
wire w0;    //: /sn:0 {0}(69,-17)(237,-17){1}
wire w3;    //: /sn:0 {0}(634,115)(661,115)(661,106)(689,106){1}
wire w104;    //: /sn:0 {0}(634,426)(670,426)(670,432)(689,432){1}
wire w111;    //: /sn:0 {0}(784,336)(794,336)(794,462)(638,462)(638,755)(727,755){1}
wire w75;    //: /sn:0 {0}(153,619)(118,619)(118,618)(111,618){1}
wire w54;    //: /sn:0 {0}(347,412)(331,412)(331,416)(253,416){1}
wire w67;    //: /sn:0 {0}(119,83)(69,83){1}
wire w90;    //: /sn:0 {0}(442,300)(457,300){1}
wire w36;    //: /sn:0 {0}(347,444)(329,444)(329,436)(253,436){1}
wire w20;    //: /sn:0 {0}(111,498)(287,498)(287,39)(351,39){1}
wire w23;    //: /sn:0 {0}(69,-27)(319,-27)(319,-9)(351,-9){1}
wire w41;    //: /sn:0 {0}(153,517)(113,517)(113,518)(111,518){1}
wire w108;    //: /sn:0 {0}(784,272)(985,272)(985,137)(1011,137){1}
wire w82;    //: /sn:0 {0}(347,396)(328,396)(328,406)(253,406){1}
wire w74;    //: /sn:0 {0}(153,609)(118,609)(118,608)(111,608){1}
wire w35;    //: /sn:0 {0}(689,-6)(649,-6)(649,-12)(634,-12){1}
wire w8;    //: /sn:0 {0}(727,643)(517,643)(517,39)(446,39){1}
wire w91;    //: /sn:0 {0}(442,316)(457,316){1}
wire w103;    //: /sn:0 {0}(634,416)(661,416)(661,416)(689,416){1}
wire w71;    //: /sn:0 {0}(347,332)(198,332)(198,578)(111,578){1}
wire w101;    //: /sn:0 {0}(634,396)(667,396)(667,384)(689,384){1}
wire w17;    //: /sn:0 {0}(634,40)(686,40)(686,42)(689,42){1}
wire w22;    //: /sn:0 {0}(351,7)(267,7)(267,478)(111,478){1}
wire w53;    //: /sn:0 {0}(1011,27)(951,27)(951,-54)(784,-54){1}
wire w84;    //: /sn:0 {0}(634,135)(672,135)(672,138)(689,138){1}
wire [3:0] w117;    //: /sn:0 {0}(#:487,260)(497,260)(497,176)(888,176)(888,82)(#:910,82){1}
wire w113;    //: /sn:0 {0}(248,132)(345,132)(345,135)(351,135){1}
wire w2;    //: /sn:0 {0}(727,739)(473,739)(473,348)(442,348){1}
wire w12;    //: /sn:0 {0}(347,364)(227,364)(227,607)(867,607)(867,659)(834,659){1}
wire w44;    //: /sn:0 {0}(69,-7)(237,-7){1}
wire w115;    //: /sn:0 {0}(248,112)(336,112)(336,103)(351,103){1}
wire w83;    //: /sn:0 {0}(634,125)(669,125)(669,122)(689,122){1}
wire w10;    //: /sn:0 {0}(834,691)(849,691){1}
wire w78;    //: /sn:0 {0}(1011,-13)(977,-13){1}
wire w27;    //: /sn:0 {0}(689,-38)(656,-38)(656,-32)(634,-32){1}
wire w52;    //: /sn:0 {0}(1011,37)(942,37)(942,-38)(784,-38){1}
wire w86;    //: /sn:0 {0}(481,245)(467,245)(467,236)(442,236){1}
wire w95;    //: /sn:0 {0}(634,298)(644,298)(644,288)(689,288){1}
wire w29;    //: /sn:0 {0}(446,23)(461,23){1}
wire w42;    //: /sn:0 {0}(69,13)(237,13){1}
wire w50;    //: /sn:0 {0}(1011,57)(920,57)(920,-6)(784,-6){1}
wire w6;    //: /sn:0 {0}(727,675)(485,675)(485,332)(442,332){1}
wire w7;    //: /sn:0 {0}(784,42)(851,42)(851,484)(697,484)(697,659)(727,659){1}
wire w93;    //: /sn:0 {0}(634,257)(654,257)(654,256)(689,256){1}
wire w112;    //: /sn:0 {0}(248,142)(335,142)(335,151)(351,151){1}
wire w46;    //: /sn:0 {0}(784,58)(861,58)(861,496)(659,496)(659,723)(727,723){1}
wire w61;    //: /sn:0 {0}(69,23)(207,23)(207,236)(347,236){1}
wire w60;    //: /sn:0 {0}(1011,97)(916,97){1}
wire w99;    //: /sn:0 {0}(689,352)(583,352)(583,565)(879,565)(879,675)(834,675){1}
wire w15;    //: /sn:0 {0}(634,30)(665,30)(665,26)(689,26){1}
wire w51;    //: /sn:0 {0}(1011,47)(929,47)(929,-22)(784,-22){1}
wire w69;    //: /sn:0 {0}(111,558)(179,558)(179,300)(347,300){1}
wire w106;    //: /sn:0 {0}(1011,117)(964,117)(964,240)(784,240){1}
wire w109;    //: /sn:0 {0}(784,288)(799,288){1}
wire w114;    //: /sn:0 {0}(248,122)(340,122)(340,119)(351,119){1}
wire w97;    //: /sn:0 {0}(634,318)(657,318)(657,320)(689,320){1}
wire w37;    //: /sn:0 {0}(689,74)(561,74)(561,573)(857,573)(857,643)(834,643){1}
wire w64;    //: /sn:0 {0}(69,53)(172,53)(172,284)(347,284){1}
wire w66;    //: /sn:0 {0}(119,73)(69,73){1}
wire w63;    //: /sn:0 {0}(347,268)(183,268)(183,43)(69,43){1}
wire w34;    //: /sn:0 {0}(1011,-3)(977,-3){1}
wire w21;    //: /sn:0 {0}(111,488)(278,488)(278,23)(351,23){1}
wire w43;    //: /sn:0 {0}(237,3)(69,3){1}
wire w76;    //: /sn:0 {0}(153,629)(118,629)(118,628)(111,628){1}
wire w87;    //: /sn:0 {0}(481,255)(458,255)(458,252)(442,252){1}
wire w102;    //: /sn:0 {0}(634,406)(676,406)(676,400)(689,400){1}
wire [3:0] w100;    //: /sn:0 {0}(#:628,35)(538,35)(538,532)(#:159,532){1}
wire w31;    //: /sn:0 {0}(446,-9)(466,-9)(466,-18)(488,-18){1}
wire w58;    //: /sn:0 {0}(153,537)(113,537)(113,538)(111,538){1}
wire w28;    //: /sn:0 {0}(689,-22)(663,-22)(663,-22)(634,-22){1}
wire w24;    //: /sn:0 {0}(69,-37)(327,-37)(327,-25)(351,-25){1}
wire [3:0] w1;    //: /sn:0 {0}(#:243,-2)(272,-2)(272,-78)(613,-78)(613,-27)(#:628,-27){1}
wire w25;    //: /sn:0 {0}(69,-47)(335,-47)(335,-41)(351,-41){1}
wire w65;    //: /sn:0 {0}(119,63)(69,63){1}
wire w98;    //: /sn:0 {0}(634,328)(644,328)(644,336)(689,336){1}
wire [3:0] w116;    //: /sn:0 {0}(#:494,-33)(559,-33)(559,-93)(963,-93)(963,2)(#:971,2){1}
wire w18;    //: /sn:0 {0}(634,50)(663,50)(663,58)(689,58){1}
wire w40;    //: /sn:0 {0}(153,527)(113,527)(113,528)(111,528){1}
wire w92;    //: /sn:0 {0}(634,247)(660,247)(660,240)(689,240){1}
wire w30;    //: /sn:0 {0}(446,7)(461,7){1}
wire w68;    //: /sn:0 {0}(119,93)(69,93){1}
wire w59;    //: /sn:0 {0}(1011,87)(916,87){1}
wire w62;    //: /sn:0 {0}(69,33)(195,33)(195,252)(347,252){1}
wire w85;    //: /sn:0 {0}(634,145)(664,145)(664,154)(689,154){1}
wire w49;    //: /sn:0 {0}(784,10)(799,10){1}
wire w57;    //: /sn:0 {0}(916,77)(1011,77){1}
wire w11;    //: /sn:0 {0}(488,-48)(467,-48)(467,-57)(446,-57){1}
wire w70;    //: /sn:0 {0}(347,316)(188,316)(188,568)(111,568){1}
wire w105;    //: /sn:0 {0}(1011,107)(952,107)(952,224)(784,224){1}
wire w72;    //: /sn:0 {0}(111,588)(209,588)(209,348)(347,348){1}
wire w88;    //: /sn:0 {0}(481,265)(462,265)(462,268)(442,268){1}
wire w94;    //: /sn:0 {0}(634,267)(644,267)(644,272)(689,272){1}
wire w13;    //: /sn:0 {0}(977,7)(1011,7){1}
wire w5;    //: /sn:0 {0}(727,691)(678,691)(678,470)(804,470)(804,320)(784,320){1}
wire w33;    //: /sn:0 {0}(488,-38)(458,-38)(458,-41)(446,-41){1}
wire w48;    //: /sn:0 {0}(784,26)(799,26){1}
wire w47;    //: /sn:0 {0}(347,428)(334,428)(334,426)(253,426){1}
wire w107;    //: /sn:0 {0}(1011,127)(975,127)(975,256)(784,256){1}
wire w9;    //: /sn:0 {0}(834,707)(849,707){1}
wire w39;    //: /sn:0 {0}(634,20)(654,20)(654,10)(689,10){1}
wire w26;    //: /sn:0 {0}(69,-57)(351,-57){1}
wire w55;    //: /sn:0 {0}(977,17)(1011,17){1}
//: enddecls

  //: IN g4 (CI) @(56,658) /sn:0 /w:[ 3 ]
  H74181 g8 (._A0(w26), ._A1(w25), ._A2(w24), ._A3(w23), ._B0(w22), ._B1(w21), ._B2(w20), ._B3(w19), .Cn(CI), .M(M), .S0(w115), .S1(w114), .S2(w113), .S3(w112), ._F0(w11), ._F1(w33), ._F2(w32), ._F3(w31), .AEB(w30), .CnP4(w29), ._G(w8), ._P(w4));   //: @(352, -73) /sz:(93, 240) /sn:0 /p:[ Li0>1 Li1>1 Li2>1 Li3>1 Li4>0 Li5>1 Li6>1 Li7>0 Li8>0 Li9>7 Li10>1 Li11>1 Li12>1 Li13>1 Ro0<1 Ro1<1 Ro2<1 Ro3<0 Ro4<0 Ro5<0 Ro6<1 Ro7<1 ]
  assign w100 = {w38, w58, w40, w41}; //: CONCAT g34  @(158,532) /sn:0 /w:[ 1 0 0 0 0 ] /dr:1 /tp:1 /drp:1
  //: OUT g3 (F) @(1050,62) /sn:0 /w:[ 1 ]
  assign {w76, w75, w74, w73, w72, w71, w70, w69, w38, w58, w40, w41, w19, w20, w21, w22} = B; //: CONCAT g13  @(106,553) /sn:0 /R:2 /w:[ 1 1 1 1 0 1 1 0 1 1 1 1 1 0 0 1 0 ] /dr:0 /tp:1 /drp:0
  //: IN g2 (OP) @(17,209) /sn:0 /w:[ 9 ]
  //: IN g1 (B) @(54,553) /sn:0 /w:[ 1 ]
  assign {w36, w47, w54, w82} = OP; //: CONCAT g16  @(248,421) /sn:0 /R:2 /w:[ 1 1 1 1 11 ] /dr:0 /tp:1 /drp:0
  assign {w68, w67, w66, w65, w64, w63, w62, w61, w42, w43, w44, w0, w23, w24, w25, w26} = A; //: CONCAT g11  @(64,18) /sn:0 /R:2 /w:[ 1 1 1 1 0 1 0 0 0 1 0 0 0 0 0 0 1 ] /dr:0 /tp:1 /drp:0
  assign {w35, w28, w27, w45} = w1; //: CONCAT g28  @(629,-27) /sn:0 /R:2 /w:[ 1 1 1 1 1 ] /dr:0 /tp:1 /drp:0
  H74181 g10 (._A0(w45), ._A1(w27), ._A2(w28), ._A3(w35), ._B0(w39), ._B1(w15), ._B2(w17), ._B3(w18), .Cn(w37), .M(M), .S0(w3), .S1(w83), .S2(w84), .S3(w85), ._F0(w53), ._F1(w52), ._F2(w51), ._F3(w50), .AEB(w49), .CnP4(w48), ._G(w7), ._P(w46));   //: @(690, -70) /sz:(93, 240) /sn:0 /p:[ Li0>0 Li1>0 Li2>0 Li3>0 Li4>1 Li5>1 Li6>1 Li7>1 Li8>0 Li9>3 Li10>1 Li11>1 Li12>1 Li13>1 Ro0<1 Ro1<1 Ro2<1 Ro3<1 Ro4<0 Ro5<0 Ro6<0 Ro7<0 ]
  assign {w98, w97, w96, w95} = w16; //: CONCAT g32  @(629,313) /sn:0 /R:2 /w:[ 0 0 0 0 0 ] /dr:0 /tp:1 /drp:0
  assign w1 = {w42, w43, w44, w0}; //: CONCAT g27  @(242,-2) /sn:0 /w:[ 0 1 0 1 1 ] /dr:1 /tp:1 /drp:1
  H74181 g19 (.S3(w36), .S2(w47), .S1(w54), .S0(w82), .M(M), .Cn(w12), ._B3(w72), ._B2(w71), ._B1(w70), ._B0(w69), ._A3(w64), ._A2(w63), ._A1(w62), ._A0(w61), ._P(w2), ._G(w6), .CnP4(w91), .AEB(w90), ._F3(w89), ._F2(w88), ._F1(w87), ._F0(w86));   //: @(348, 220) /sz:(93, 240) /sn:0 /p:[ Li0>0 Li1>0 Li2>0 Li3>0 Li4>11 Li5>0 Li6>1 Li7>0 Li8>0 Li9>1 Li10>1 Li11>0 Li12>1 Li13>1 Ro0<1 Ro1<1 Ro2<0 Ro3<0 Ro4<1 Ro5<1 Ro6<1 Ro7<1 ]
  //: IN g6 (M) @(12,183) /sn:0 /w:[ 9 ]
  H74182 g7 (._G0(w8), ._G1(w7), ._G2(w6), ._G3(w5), ._P0(w4), ._P1(w46), ._P2(w2), ._P3(w111), .Cn(CI), .CnPx(w37), .CnPy(w12), .CnPz(w99), ._G(w10), ._P(w9));   //: @(728, 627) /sz:(105, 160) /sn:0 /p:[ Li0>0 Li1>1 Li2>0 Li3>0 Li4>0 Li5>1 Li6>0 Li7>1 Li8>5 Ro0<1 Ro1<1 Ro2<1 Ro3<0 Ro4<0 ]
  //: joint g9 (CI) @(325, 657) /w:[ -1 1 2 4 ]
  //: joint g15 (OP) @(218, 209) /w:[ 5 6 8 10 ]
  assign w16 = {w76, w75, w74, w73}; //: CONCAT g31  @(158,614) /sn:0 /w:[ 1 0 0 0 0 ] /dr:1 /tp:1 /drp:1
  H74181 g20 (.S3(w104), .S2(w103), .S1(w102), .S0(w101), .M(M), .Cn(w99), ._B3(w98), ._B2(w97), ._B1(w96), ._B0(w95), ._A3(w94), ._A2(w93), ._A1(w92), ._A0(w81), ._P(w111), ._G(w5), .CnP4(CO), .AEB(w109), ._F3(w108), ._F2(w107), ._F1(w106), ._F0(w105));   //: @(690, 208) /sz:(93, 240) /sn:0 /p:[ Li0>1 Li1>1 Li2>1 Li3>1 Li4>0 Li5>0 Li6>1 Li7>1 Li8>1 Li9>1 Li10>1 Li11>1 Li12>1 Li13>1 Ro0<0 Ro1<1 Ro2<1 Ro3<0 Ro4<0 Ro5<1 Ro6<1 Ro7<1 ]
  assign {w55, w13, w34, w78} = w116; //: CONCAT g25  @(972,2) /sn:0 /R:2 /w:[ 0 0 1 1 1 ] /dr:0 /tp:1 /drp:0
  assign {w85, w84, w83, w3} = OP; //: CONCAT g17  @(629,130) /sn:0 /R:2 /w:[ 0 0 0 0 3 ] /dr:0 /tp:1 /drp:0
  assign w14 = {w68, w67, w66, w65}; //: CONCAT g29  @(124,78) /sn:0 /w:[ 0 0 0 0 0 ] /dr:1 /tp:1 /drp:1
  assign {w112, w113, w114, w115} = OP; //: CONCAT g14  @(243,127) /sn:0 /R:2 /w:[ 0 0 0 0 7 ] /dr:0 /tp:1 /drp:0
  //: OUT g5 (CO) @(991,307) /sn:0 /w:[ 0 ]
  assign w117 = {w89, w88, w87, w86}; //: CONCAT g24  @(486,260) /sn:0 /w:[ 0 0 0 0 0 ] /dr:1 /tp:1 /drp:1
  assign {w104, w103, w102, w101} = OP; //: CONCAT g21  @(629,411) /sn:0 /R:2 /w:[ 0 0 0 0 0 ] /dr:0 /tp:1 /drp:0
  assign {w60, w59, w57, w56} = w117; //: CONCAT g23  @(911,82) /sn:0 /R:2 /w:[ 1 1 0 0 1 ] /dr:0 /tp:1 /drp:0
  assign w116 = {w31, w32, w33, w11}; //: CONCAT g35  @(493,-33) /sn:0 /w:[ 0 1 0 0 0 ] /dr:1 /tp:1 /drp:1
  //: joint g22 (OP) @(595, 209) /w:[ -1 2 4 1 ]
  //: joint g26 (M) @(571, 183) /w:[ -1 2 4 1 ]
  //: IN g0 (A) @(12,18) /sn:0 /w:[ 0 ]
  //: joint g12 (M) @(312, 183) /w:[ 5 6 8 10 ]
  assign F = {w108, w107, w106, w105, w60, w59, w57, w56, w50, w51, w52, w53, w55, w13, w34, w78}; //: CONCAT g18  @(1016,62) /sn:0 /w:[ 0 1 0 0 0 0 0 1 1 0 0 0 0 1 1 0 0 ] /dr:1 /tp:1 /drp:1
  assign {w18, w17, w15, w39} = w100; //: CONCAT g33  @(629,35) /sn:0 /R:2 /w:[ 0 0 0 0 0 ] /dr:0 /tp:1 /drp:0
  assign {w94, w93, w92, w81} = w14; //: CONCAT g30  @(629,252) /sn:0 /R:2 /w:[ 0 0 0 0 1 ] /dr:0 /tp:1 /drp:0

endmodule
//: /netlistEnd


//: version "2.0-b10"
//: property encoding = "iso8859-1"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "stdlogic.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"
//: require "74xx"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg [15:0] A_NET;    //: {0}(#:50:157,129)(206,129)(206,167)(249,167){1}
reg w0;    //: /sn:0 {0}(130,199)(249,199){1}
reg [3:0] w18;    //: /sn:0 {0}(#:154,239)(202,239)(202,215)(249,215){1}
wire [15:0] w4;    //: /sn:0 {0}(413,183)(355,183){1}
wire [15:0] w2;    //: /sn:0 {0}(#:234,183)(249,183){1}
wire w5;    //: /sn:0 {0}(387,167)(355,167){1}
//: enddecls

  //: SWITCH M (w0) @(113,199) /w:[ 0 ] /st:1 /dn:1
  //: LED g1 (w5) @(394,167) /sn:0 /R:3 /w:[ 0 ] /type:0
  //: DIP A (A_NET) @(119,129) /R:1 /w:[ 0 ] /st:2 /dn:1
  //: LED g6 (w4) @(420,183) /sn:0 /R:3 /w:[ 0 ] /type:2
  //: DIP OP (w18) @(116,239) /R:1 /w:[ 0 ] /st:0 /dn:1
  ALU16_74181 g0 (.A(A_NET), .B(w2), .M(w0), .S(w18), .C(w5), .F(w4));   //: @(250, 151) /sz:(104, 80) /sn:0 /p:[ Li0>1 Li1>1 Li2>1 Li3>1 Ro0<1 Ro1<1 ]

endmodule
//: /netlistEnd

//: /netlistBegin ALU16_74181
module ALU16_74181(F, S, M, B, C, A);
//: interface  /sz:(104, 80) /bd:[ Li0>S[3:0](64/80) Li1>M(48/80) Li2>B[15:0](32/80) Li3>A[15:0](16/80) Ro0<F[15:0](32/80) Ro1<C(16/80) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input M;    //: {0}(413,197)(326,197)(326,190)(33,190)(33,366){1}
//: {2}(35,368)(51,368){3}
//: {4}(53,366)(53,199)(119,199){5}
//: {6}(53,370)(53,563)(119,563){7}
//: {8}(31,368)(21,368)(21,367)(99:-194,367){9}
//: {10}(33,370)(33,557)(453,557){11}
input [15:0] B;    //: /sn:0 {0}(#:-226,481)(-211,481){1}
output [15:0] F;    //: /sn:0 {0}(771,253)(#:704,253){1}
input [15:0] A;    //: {0}(#:80:-175,129)(#:58:-101,129){1}
output C;    //: /sn:0 {0}(787,463)(731,463)(731,493)(548,493){1}
supply0 w2;    //: /sn:0 {0}(62,163)(62,183)(119,183){1}
input [3:0] S;    //: {0}(#:70:-216,290)(#:-139,290){1}
wire w32;    //: /sn:0 {0}(-95,164)(-3,164)(-3,467)(119,467){1}
wire w6;    //: /sn:0 {0}(119,167)(104,167){1}
wire w73;    //: /sn:0 {0}(453,509)(433,509){1}
wire w45;    //: /sn:0 {0}(453,605)(363,605)(363,390)(167,390)(167,331){1}
//: {2}(169,329)(359,329)(359,245)(413,245){3}
//: {4}(165,329)(48,329)(48,297){5}
//: {6}(48,293)(48,247)(119,247){7}
//: {8}(46,295)(-74,295){9}
//: {10}(-78,295)(-133,295){11}
//: {12}(-76,297)(-76,611)(119,611){13}
wire w93;    //: /sn:0 {0}(508,85)(622,85)(622,238)(698,238){1}
wire w96;    //: /sn:0 {0}(214,435)(337,435)(337,375)(581,375)(581,268)(698,268){1}
wire w7;    //: /sn:0 {0}(119,151)(104,151){1}
wire w46;    //: /sn:0 {0}(413,229)(350,229)(350,319)(203,319){1}
//: {2}(199,319)(39,319)(39,287){3}
//: {4}(39,283)(39,231)(119,231){5}
//: {6}(37,285)(-64,285){7}
//: {8}(-68,285)(-133,285){9}
//: {10}(-66,287)(-66,595)(119,595){11}
//: {12}(201,321)(201,379)(371,379)(371,589)(453,589){13}
wire w99;    //: /sn:0 {0}(698,298)(614,298)(614,413)(548,413){1}
wire w61;    //: /sn:0 {0}(508,117)(523,117){1}
wire w60;    //: /sn:0 {0}(119,547)(109,547)(109,532)(188,532)(188,357)(545,357)(545,133)(508,133){1}
wire w56;    //: /sn:0 {0}(-95,104)(45,104)(45,-51)(384,-51)(384,69)(413,69){1}
wire w16;    //: /sn:0 {0}(214,135)(351,135)(351,181)(413,181){1}
wire w14;    //: /sn:0 {0}(214,167)(229,167){1}
wire w81;    //: /sn:0 {0}(548,509)(563,509){1}
wire w19;    //: /sn:0 {0}(214,87)(257,87)(257,19)(662,19)(662,198)(698,198){1}
wire w15;    //: /sn:0 {0}(214,151)(229,151){1}
wire w38;    //: /sn:0 {0}(214,499)(398,499)(398,541)(453,541){1}
wire w51;    //: /sn:0 {0}(413,149)(398,149){1}
wire w0;    //: /sn:0 {0}(453,621)(335,621)(335,397)(148,397)(148,340){1}
//: {2}(150,338)(370,338)(370,261)(413,261){3}
//: {4}(146,338)(57,338)(57,307){5}
//: {6}(57,303)(57,263)(119,263){7}
//: {8}(55,305)(-89,305){9}
//: {10}(-93,305)(-133,305){11}
//: {12}(-91,307)(-91,627)(119,627){13}
wire w97;    //: /sn:0 {0}(214,451)(348,451)(348,386)(591,386)(591,278)(698,278){1}
wire w64;    //: /sn:0 {0}(508,69)(633,69)(633,228)(698,228){1}
wire w37;    //: /sn:0 {0}(214,515)(229,515){1}
wire w34;    //: /sn:0 {0}(-95,144)(12,144)(12,435)(119,435){1}
wire w76;    //: /sn:0 {0}(453,461)(430,461)(430,692)(63,692)(63,204)(-95,204){1}
wire w75;    //: /sn:0 {0}(453,477)(438,477){1}
wire w102;    //: /sn:0 {0}(548,461)(649,461)(649,328)(698,328){1}
wire w43;    //: /sn:0 {0}(214,419)(328,419)(328,366)(572,366)(572,258)(698,258){1}
wire w21;    //: /sn:0 {0}(214,55)(235,55)(235,-5)(683,-5)(683,178)(698,178){1}
wire w54;    //: /sn:0 {0}(-95,124)(69,124)(69,-27)(364,-27)(364,101)(413,101){1}
wire w100;    //: /sn:0 {0}(548,429)(625,429)(625,308)(698,308){1}
wire w58;    //: /sn:0 {0}(508,165)(523,165){1}
wire w31;    //: /sn:0 {0}(119,483)(104,483){1}
wire w90;    //: /sn:0 {0}(214,103)(358,103)(358,31)(651,31)(651,208)(698,208){1}
wire w28;    //: /sn:0 {0}(119,531)(104,531){1}
wire w36;    //: /sn:0 {0}(214,531)(229,531){1}
wire w20;    //: /sn:0 {0}(214,71)(246,71)(246,7)(673,7)(673,188)(698,188){1}
wire w1;    //: /sn:0 {0}(453,573)(381,573)(381,351)(229,351)(229,313){1}
//: {2}(231,311)(345,311)(345,213)(413,213){3}
//: {4}(227,311)(29,311)(29,277){5}
//: {6}(29,273)(29,215)(119,215){7}
//: {8}(27,275)(-55,275){9}
//: {10}(-59,275)(-133,275){11}
//: {12}(-57,277)(-57,579)(119,579){13}
wire w74;    //: /sn:0 {0}(453,493)(438,493){1}
wire w65;    //: /sn:0 {0}(508,53)(642,53)(642,218)(698,218){1}
wire w98;    //: /sn:0 {0}(698,288)(601,288)(601,395)(358,395)(358,467)(214,467){1}
wire w35;    //: /sn:0 {0}(-95,134)(22,134)(22,419)(119,419){1}
wire w8;    //: /sn:0 {0}(119,135)(104,135){1}
wire w101;    //: /sn:0 {0}(698,318)(635,318)(635,445)(548,445){1}
wire w30;    //: /sn:0 {0}(119,499)(104,499){1}
wire w17;    //: /sn:0 {0}(214,119)(229,119){1}
wire w53;    //: /sn:0 {0}(413,117)(398,117){1}
wire w59;    //: /sn:0 {0}(508,149)(523,149){1}
wire w62;    //: /sn:0 {0}(508,101)(613,101)(613,248)(698,248){1}
wire w57;    //: /sn:0 {0}(-95,94)(33,94)(33,-63)(394,-63)(394,53)(413,53){1}
wire w12;    //: /sn:0 {0}(-95,64)(104,64)(104,71)(119,71){1}
wire w11;    //: /sn:0 {0}(-95,74)(94,74)(94,87)(119,87){1}
wire w77;    //: /sn:0 {0}(453,445)(420,445)(420,683)(74,683)(74,194)(-95,194){1}
wire w83;    //: /sn:0 {0}(548,477)(563,477){1}
wire w78;    //: /sn:0 {0}(-95,184)(82,184)(82,674)(412,674)(412,429)(453,429){1}
wire w10;    //: /sn:0 {0}(-95,84)(87,84)(87,103)(119,103){1}
wire w72;    //: /sn:0 {0}(453,525)(438,525){1}
wire w13;    //: /sn:0 {0}(-95,54)(104,54)(104,55)(119,55){1}
wire w52;    //: /sn:0 {0}(413,133)(398,133){1}
wire w33;    //: /sn:0 {0}(-95,154)(4,154)(4,451)(119,451){1}
wire w80;    //: /sn:0 {0}(548,525)(602,525){1}
wire w29;    //: /sn:0 {0}(119,515)(104,515){1}
wire w79;    //: /sn:0 {0}(-95,174)(90,174)(90,666)(403,666)(403,413)(453,413){1}
wire w50;    //: /sn:0 {0}(413,165)(398,165){1}
wire w9;    //: /sn:0 {0}(119,119)(104,119){1}
wire w55;    //: /sn:0 {0}(-95,114)(57,114)(57,-39)(374,-39)(374,85)(413,85){1}
wire w39;    //: /sn:0 {0}(214,483)(229,483){1}
//: enddecls

  //: OUT g4 (F) @(768,253) /sn:0 /w:[ 0 ]
  //: joint g8 (w1) @(-57, 275) /w:[ 9 -1 10 12 ]
  //: IN g3 (S) @(-218,290) /sn:0 /w:[ 0 ]
  //: joint g13 (w46) @(39, 285) /w:[ -1 4 6 3 ]
  //: IN g2 (M) @(-196,367) /sn:0 /w:[ 9 ]
  //: IN g1 (B) @(-228,481) /sn:0 /w:[ 0 ]
  H74181 g11 (._A0(w35), ._A1(w34), ._A2(w33), ._A3(w32), ._B0(w31), ._B1(w30), ._B2(w29), ._B3(w28), .Cn(w60), .M(M), .S0(w1), .S1(w46), .S2(w45), .S3(w0), ._F0(w43), ._F1(w96), ._F2(w97), ._F3(w98), .AEB(w39), .CnP4(w38), ._G(w37), ._P(w36));   //: @(120, 403) /sz:(93, 240) /sn:0 /p:[ Li0>1 Li1>1 Li2>1 Li3>1 Li4>0 Li5>0 Li6>0 Li7>0 Li8>0 Li9>7 Li10>13 Li11>11 Li12>13 Li13>13 Ro0<0 Ro1<0 Ro2<0 Ro3<1 Ro4<0 Ro5<0 Ro6<0 Ro7<0 ]
  //: joint g16 (w1) @(229, 311) /w:[ 2 -1 4 1 ]
  H74181 g10 (._A0(w57), ._A1(w56), ._A2(w55), ._A3(w54), ._B0(w53), ._B1(w52), ._B2(w51), ._B3(w50), .Cn(w16), .M(M), .S0(w1), .S1(w46), .S2(w45), .S3(w0), ._F0(w65), ._F1(w64), ._F2(w93), ._F3(w62), .AEB(w61), .CnP4(w60), ._G(w59), ._P(w58));   //: @(414, 37) /sz:(93, 240) /sn:0 /p:[ Li0>1 Li1>1 Li2>1 Li3>1 Li4>0 Li5>0 Li6>0 Li7>0 Li8>1 Li9>0 Li10>3 Li11>0 Li12>3 Li13>3 Ro0<0 Ro1<0 Ro2<0 Ro3<0 Ro4<0 Ro5<1 Ro6<0 Ro7<0 ]
  //: joint g28 (w45) @(167, 329) /w:[ 2 -1 4 1 ]
  //: joint g19 (w0) @(148, 338) /w:[ 2 -1 4 1 ]
  H74181 g9 (._A0(w79), ._A1(w78), ._A2(w77), ._A3(w76), ._B0(w75), ._B1(w74), ._B2(w73), ._B3(w72), .Cn(w38), .M(M), .S0(w1), .S1(w46), .S2(w45), .S3(w0), ._F0(w99), ._F1(w100), ._F2(w101), ._F3(w102), .AEB(w83), .CnP4(C), ._G(w81), ._P(w80));   //: @(454, 397) /sz:(93, 240) /sn:0 /p:[ Li0>1 Li1>1 Li2>0 Li3>0 Li4>0 Li5>0 Li6>0 Li7>0 Li8>1 Li9>11 Li10>0 Li11>13 Li12>0 Li13>0 Ro0<1 Ro1<0 Ro2<1 Ro3<0 Ro4<0 Ro5<1 Ro6<0 Ro7<0 ]
  //: joint g7 (w0) @(-91, 305) /w:[ 9 -1 10 12 ]
  //: joint g15 (w46) @(-66, 285) /w:[ 7 -1 8 10 ]
  //: GROUND g20 (w2) @(62,157) /sn:0 /R:2 /w:[ 0 ]
  assign {w76, w77, w78, w79, w32, w33, w34, w35, w54, w55, w56, w57, w10, w11, w12, w13} = A; //: CONCAT g17  @(-100,129) /sn:0 /R:2 /w:[ 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 ] /dr:0 /tp:1 /drp:0
  H74181 g29 (._A0(w13), ._A1(w12), ._A2(w11), ._A3(w10), ._B0(w9), ._B1(w8), ._B2(w7), ._B3(w6), .Cn(w2), .M(M), .S0(w1), .S1(w46), .S2(w45), .S3(w0), ._F0(w21), ._F1(w20), ._F2(w19), ._F3(w90), .AEB(w17), .CnP4(w16), ._G(w15), ._P(w14));   //: @(120, 39) /sz:(93, 240) /sn:0 /p:[ Li0>1 Li1>1 Li2>1 Li3>1 Li4>0 Li5>0 Li6>0 Li7>0 Li8>1 Li9>5 Li10>7 Li11>5 Li12>7 Li13>7 Ro0<0 Ro1<0 Ro2<0 Ro3<0 Ro4<0 Ro5<0 Ro6<0 Ro7<0 ]
  //: OUT g5 (C) @(784,463) /sn:0 /w:[ 0 ]
  assign {w0, w45, w46, w1} = S; //: CONCAT g14  @(-138,290) /sn:0 /R:2 /w:[ 11 11 9 11 1 ] /dr:0 /tp:1 /drp:0
  //: joint g21 (w46) @(201, 319) /w:[ 1 -1 2 12 ]
  //: joint g24 (M) @(33, 368) /w:[ 2 1 8 10 ]
  assign F = {w102, w101, w100, w99, w98, w97, w96, w43, w62, w93, w64, w65, w90, w19, w20, w21}; //: CONCAT g23  @(703,253) /sn:0 /w:[ 1 1 0 1 0 0 1 1 1 1 1 1 1 1 1 1 1 ] /dr:1 /tp:1 /drp:1
  //: IN g0 (A) @(-177,129) /sn:0 /w:[ 0 ]
  //: joint g22 (w45) @(48, 295) /w:[ -1 6 8 5 ]
  //: joint g26 (M) @(53, 368) /w:[ -1 4 3 6 ]
  //: joint g12 (w45) @(-76, 295) /w:[ 9 -1 10 12 ]
  //: joint g18 (w0) @(57, 305) /w:[ -1 6 8 5 ]
  //: joint g30 (w1) @(29, 275) /w:[ -1 6 8 5 ]

endmodule
//: /netlistEnd


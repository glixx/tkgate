//: version "2.1"
//: property encoding = "utf-8"
//: property locale = "uk"
//: property prefix = "_GG"
//: property title = "Combinational Simulation"
//: property useExtBars = 0
//: property showSwitchNets = 0
//: property discardChanges = 1
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin PAGE1
module PAGE1;    //: root_module
//: enddecls

  //: comment g13 @(10,10) /anc:1
  //: /line:"<h3>Combinational Circuit Simulation</h3>"
  //: /line:""
  //: /line:"TkGate uses a Verilog-based discrete event simulator to simulate your circuit description. In this"
  //: /line:"chapter the basics needed to simulate a combinational circuit will be presented."
  //: /end
  //: comment g0 @(191,165) /sn:0 /anc:1
  //: /line:"<img src=simulate.gif>"
  //: /end
  //: comment g12 @(10,410) /sn:0 /R:14 /anc:1
  //: /line:"<tutorial-navigation byfile=1>"
  //: /end

endmodule
//: /netlistEnd


//: version "2.1-a2"
//: property encoding = "utf-8"
//: property locale = "it"
//: property prefix = "_GG"
//: property title = "Sequential Simulation"
//: property useExtBars = 0
//: property showSwitchNets = 0
//: property discardChanges = 1
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin PAGE1
module PAGE1;    //: root_module
//: enddecls

  //: comment g13 @(14,12) /anc:1
  //: /line:"<h3>Sequential Simulation</h3>"
  //: /line:""
  //: /line:"This chapter builds on the previous chapter about simulating combinational circuits and introduces"
  //: /line:"simulator features that are useful for simulating sequential circuits."
  //: /end
  //: comment g1 @(10,410) /sn:0 /R:14 /anc:1
  //: /line:"<tutorial-navigation byfile=1>"
  //: /end
  //: comment g10 @(208,188) /sn:0 /anc:1
  //: /line:"<img src=simulate.gif>"
  //: /end

endmodule
//: /netlistEnd


//: version "2.0-b10"
//: property encoding = "iso8859-1"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "74 series standart logic circuits"
//: property showSwitchNets = 0
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg w45;    //: /sn:0 {0}(822,167)(761,167)(761,135)(647,135){1}
reg w166;    //: /sn:0 {0}(1008,495)(1067,495)(1067,571)(1089,571){1}
reg w134;    //: /sn:0 {0}(51,1021)(77,1021)(77,1084){1}
//: {2}(79,1086)(317,1086){3}
//: {4}(77,1088)(77,1240)(317,1240){5}
reg w14;    //: /sn:0 {0}(634,658)(658,658)(658,644)(718,644){1}
reg w89;    //: /sn:0 {0}(637,1049)(705,1049)(705,964)(735,964){1}
reg w4;    //: /sn:0 {0}(773,705)(773,768)(721,768){1}
reg w38;    //: /sn:0 {0}(319,1529)(252,1529){1}
//: {2}(250,1527)(250,1339){3}
//: {4}(252,1337)(316,1337){5}
//: {6}(250,1335)(250,840){7}
//: {8}(252,838)(316,838){9}
//: {10}(250,836)(250,667){11}
//: {12}(252,665)(314,665){13}
//: {14}(250,663)(250,512){15}
//: {16}(252,510)(312,510){17}
//: {18}(250,508)(250,390){19}
//: {20}(252,388)(309,388){21}
//: {22}(250,386)(250,237){23}
//: {24}(252,235)(310,235){25}
//: {26}(250,233)(250,84){27}
//: {28}(252,82)(310,82){29}
//: {30}(248,82)(106,82)(106,134)(63,134){31}
//: {32}(250,1531)(250,1682){33}
//: {34}(252,1684)(317,1684){35}
//: {36}(250,1686)(250,1881){37}
//: {38}(252,1883)(319,1883){39}
//: {40}(250,1885)(250,2035)(319,2035){41}
reg w152;    //: /sn:0 {0}(1085,307)(1048,307)(1048,422)(980,422){1}
reg w151;    //: /sn:0 {0}(1085,195)(1003,195)(1003,186)(981,186){1}
reg w0;    //: /sn:0 {0}(316,854)(223,854){1}
//: {2}(221,852)(221,683){3}
//: {4}(223,681)(314,681){5}
//: {6}(221,679)(221,544){7}
//: {8}(223,542)(312,542){9}
//: {10}(221,540)(221,269){11}
//: {12}(223,267)(310,267){13}
//: {14}(221,265)(221,116){15}
//: {16}(223,114)(310,114){17}
//: {18}(219,114)(129,114)(129,231)(63,231){19}
//: {20}(221,856)(221,1004){21}
//: {22}(223,1006)(317,1006){23}
//: {24}(221,1008)(221,1157){25}
//: {26}(223,1159)(233,1159)(233,1160)(317,1160){27}
//: {28}(221,1161)(221,1351){29}
//: {30}(223,1353)(316,1353){31}
//: {32}(221,1355)(221,1559){33}
//: {34}(223,1561)(319,1561){35}
//: {36}(221,1563)(221,1913){37}
//: {38}(223,1915)(319,1915){39}
//: {40}(221,1917)(221,2067)(319,2067){41}
reg w3;    //: /sn:0 {0}(310,315)(183,315){1}
//: {2}(181,313)(181,164){3}
//: {4}(183,162)(310,162){5}
//: {6}(179,162)(167,162)(167,354)(63,354){7}
//: {8}(181,317)(181,588){9}
//: {10}(183,590)(312,590){11}
//: {12}(181,592)(181,1607){13}
//: {14}(183,1609)(319,1609){15}
//: {16}(181,1611)(181,1787)(180,1787)(180,1961){17}
//: {18}(182,1963)(319,1963){19}
//: {20}(180,1965)(180,2115)(319,2115){21}
reg w120;    //: /sn:0 {0}(734,1705)(753,1705)(753,1666){1}
reg w171;    //: /sn:0 {0}(1008,673)(1027,673)(1027,635)(1089,635){1}
reg w168;    //: /sn:0 {0}(1089,619)(1008,619){1}
reg w133;    //: /sn:0 {0}(51,976)(91,976)(91,1068){1}
//: {2}(93,1070)(317,1070){3}
//: {4}(91,1072)(91,1224)(317,1224){5}
reg w111;    //: /sn:0 {0}(621,1537)(659,1537)(659,1537)(700,1537){1}
reg w90;    //: /sn:0 {0}(621,1622)(660,1622)(660,1585)(700,1585){1}
reg w167;    //: /sn:0 {0}(1008,578)(1033,578)(1033,603)(1089,603){1}
reg w36;    //: /sn:0 {0}(316,806)(282,806){1}
//: {2}(280,804)(280,635){3}
//: {4}(282,633)(314,633){5}
//: {6}(280,631)(280,480){7}
//: {8}(282,478)(312,478){9}
//: {10}(280,476)(280,358){11}
//: {12}(282,356)(309,356){13}
//: {14}(280,354)(280,205){15}
//: {16}(282,203)(310,203){17}
//: {18}(280,201)(280,52){19}
//: {20}(282,50)(310,50){21}
//: {22}(278,50)(63,50){23}
//: {24}(280,808)(280,972){25}
//: {26}(282,974)(317,974){27}
//: {28}(280,976)(280,1126){29}
//: {30}(282,1128)(317,1128){31}
//: {32}(280,1130)(280,1303){33}
//: {34}(282,1305)(316,1305){35}
//: {36}(280,1307)(280,1495){37}
//: {38}(282,1497)(319,1497){39}
//: {40}(280,1499)(280,1650){41}
//: {42}(282,1652)(317,1652){43}
//: {44}(280,1654)(280,1849){45}
//: {46}(282,1851)(319,1851){47}
//: {48}(280,1853)(280,2003)(319,2003){49}
reg w41;    //: /sn:0 {0}(66,420)(309,420){1}
reg w108;    //: /sn:0 {0}(619,1300)(635,1300)(635,1328)(693,1328){1}
reg w126;    //: /sn:0 {0}(1007,841)(1074,841)(1074,699)(1089,699){1}
reg w91;    //: /sn:0 {0}(729,1495)(755,1495)(755,1425){1}
reg w144;    //: /sn:0 {0}(981,18)(1067,18)(1067,115)(1085,115){1}
reg w84;    //: /sn:0 {0}(637,867)(720,867)(720,884)(735,884){1}
reg w172;    //: /sn:0 {0}(1008,714)(1039,714)(1039,651)(1089,651){1}
reg w2;    //: /sn:0 {0}(316,1385)(197,1385){1}
//: {2}(195,1383)(195,889){3}
//: {4}(197,887)(207,887)(207,886)(316,886){5}
//: {6}(195,885)(195,715){7}
//: {8}(197,713)(314,713){9}
//: {10}(195,711)(195,576){11}
//: {12}(197,574)(312,574){13}
//: {14}(195,572)(195,301){15}
//: {16}(197,299)(310,299){17}
//: {18}(195,297)(195,148){19}
//: {20}(197,146)(310,146){21}
//: {22}(193,146)(154,146)(154,313)(63,313){23}
//: {24}(195,1387)(195,1591){25}
//: {26}(197,1593)(319,1593){27}
//: {28}(195,1595)(195,1945){29}
//: {30}(197,1947)(319,1947){31}
//: {32}(195,1949)(195,2099)(319,2099){33}
reg w12;    //: /sn:0 {0}(316,918)(154,918){1}
//: {2}(152,916)(152,747){3}
//: {4}(154,745)(314,745){5}
//: {6}(150,745)(78,745)(78,772)(55,772){7}
//: {8}(152,920)(152,1052){9}
//: {10}(154,1054)(317,1054){11}
//: {12}(152,1056)(152,1206){13}
//: {14}(154,1208)(317,1208){15}
//: {16}(152,1210)(152,1417)(316,1417){17}
reg w44;    //: /sn:0 {0}(822,151)(790,151)(790,91)(648,91){1}
reg w86;    //: /sn:0 {0}(637,941)(664,941)(664,916)(735,916){1}
reg w155;    //: /sn:0 {0}(1085,291)(1041,291)(1041,390)(980,390){1}
reg w147;    //: /sn:0 {0}(981,114)(1026,114)(1026,163)(1085,163){1}
reg w50;    //: /sn:0 {0}(648,368)(727,368)(727,247)(822,247){1}
reg w6;    //: /sn:0 {0}(635,690)(673,690)(673,660)(718,660){1}
reg w7;    //: /sn:0 {0}(316,902)(168,902){1}
//: {2}(166,900)(166,731){3}
//: {4}(168,729)(314,729){5}
//: {6}(164,729)(56,729){7}
//: {8}(166,904)(166,1008)(166,1008)(166,1036){9}
//: {10}(168,1038)(317,1038){11}
//: {12}(166,1040)(166,1190){13}
//: {14}(168,1192)(317,1192){15}
//: {16}(166,1194)(166,1401)(316,1401){17}
reg w93;    //: /sn:0 {0}(693,1360)(650,1360)(650,1399)(610,1399){1}
reg w61;    //: /sn:0 {0}(319,2131)(148,2131){1}
reg w46;    //: /sn:0 {0}(822,183)(648,183){1}
reg w99;    //: /sn:0 {0}(693,1392)(677,1392)(677,1466)(610,1466){1}
reg w153;    //: /sn:0 {0}(980,455)(1055,455)(1055,323)(1085,323){1}
reg w15;    //: /sn:0 {0}(634,604)(665,604)(665,628)(718,628){1}
reg w106;    //: /sn:0 {0}(693,1296)(653,1296)(653,1241)(619,1241){1}
reg w109;    //: /sn:0 {0}(621,1593)(652,1593)(652,1569)(700,1569){1}
reg w37;    //: /sn:0 {0}(316,822)(268,822){1}
//: {2}(266,820)(266,651){3}
//: {4}(268,649)(314,649){5}
//: {6}(266,647)(266,496){7}
//: {8}(268,494)(312,494){9}
//: {10}(266,492)(266,374){11}
//: {12}(268,372)(309,372){13}
//: {14}(266,370)(266,221){15}
//: {16}(268,219)(310,219){17}
//: {18}(266,217)(266,68){19}
//: {20}(268,66)(310,66){21}
//: {22}(264,66)(92,66)(92,91)(63,91){23}
//: {24}(266,824)(266,988){25}
//: {26}(268,990)(317,990){27}
//: {28}(266,992)(266,1141){29}
//: {30}(268,1143)(278,1143)(278,1144)(317,1144){31}
//: {32}(266,1145)(266,1319){33}
//: {34}(268,1321)(316,1321){35}
//: {36}(266,1323)(266,1511){37}
//: {38}(268,1513)(319,1513){39}
//: {40}(266,1515)(266,1666){41}
//: {42}(268,1668)(317,1668){43}
//: {44}(266,1670)(266,1865){45}
//: {46}(268,1867)(319,1867){47}
//: {48}(266,1869)(266,2019)(319,2019){49}
reg w159;    //: /sn:0 {0}(1089,587)(1051,587)(1051,536)(1008,536){1}
reg w63;    //: /sn:0 {0}(621,1663)(666,1663)(666,1601)(700,1601){1}
reg w87;    //: /sn:0 {0}(637,977)(674,977)(674,932)(735,932){1}
reg w43;    //: /sn:0 {0}(649,44)(807,44)(807,135)(822,135){1}
reg w170;    //: /sn:0 {0}(1089,683)(1060,683)(1060,797)(1008,797){1}
reg w58;    //: /sn:0 {0}(635,543)(700,543)(700,596)(718,596){1}
reg w169;    //: /sn:0 {0}(1008,756)(1048,756)(1048,667)(1089,667){1}
reg w28;    //: /sn:0 {0}(981,296)(1026,296)(1026,243)(1085,243){1}
reg w24;    //: /sn:0 {0}(634,574)(681,574)(681,612)(718,612){1}
reg w1;    //: /sn:0 {0}(316,870)(211,870){1}
//: {2}(209,868)(209,699){3}
//: {4}(211,697)(314,697){5}
//: {6}(209,695)(209,560){7}
//: {8}(211,558)(312,558){9}
//: {10}(209,556)(209,285){11}
//: {12}(211,283)(310,283){13}
//: {14}(209,281)(209,132){15}
//: {16}(211,130)(310,130){17}
//: {18}(207,130)(142,130)(142,272)(63,272){19}
//: {20}(209,872)(209,1020){21}
//: {22}(211,1022)(317,1022){23}
//: {24}(209,1024)(209,1173){25}
//: {26}(211,1175)(221,1175)(221,1176)(317,1176){27}
//: {28}(209,1177)(209,1366){29}
//: {30}(211,1368)(221,1368)(221,1369)(316,1369){31}
//: {32}(209,1370)(209,1575){33}
//: {34}(211,1577)(319,1577){35}
//: {36}(209,1579)(209,1929){37}
//: {38}(211,1931)(319,1931){39}
//: {40}(209,1933)(209,2083)(319,2083){41}
reg w154;    //: /sn:0 {0}(980,359)(1034,359)(1034,275)(1085,275){1}
reg w121;    //: /sn:0 {0}(700,1553)(644,1553)(644,1565)(621,1565){1}
reg w40;    //: /sn:0 {0}(66,460)(76,460)(76,436)(309,436){1}
reg w92;    //: /sn:0 {0}(693,1344)(625,1344)(625,1366)(610,1366){1}
reg w149;    //: /sn:0 {0}(981,155)(1021,155)(1021,179)(1085,179){1}
reg w146;    //: /sn:0 {0}(981,81)(1040,81)(1040,147)(1085,147){1}
reg w59;    //: /sn:0 {0}(148,2162)(304,2162)(304,2147)(319,2147){1}
reg w62;    //: /sn:0 {0}(981,324)(1030,324)(1030,259)(1085,259){1}
reg w85;    //: /sn:0 {0}(735,900)(652,900)(652,905)(637,905){1}
reg w49;    //: /sn:0 {0}(648,322)(698,322)(698,231)(822,231){1}
reg w150;    //: /sn:0 {0}(1085,211)(993,211)(993,218)(981,218){1}
reg w148;    //: /sn:0 {0}(981,251)(1019,251)(1019,227)(1085,227){1}
reg w105;    //: /sn:0 {0}(693,1280)(674,1280)(674,1212)(619,1212){1}
reg w110;    //: /sn:0 {0}(621,1688)(674,1688)(674,1617)(700,1617){1}
reg w88;    //: /sn:0 {0}(637,1013)(687,1013)(687,948)(735,948){1}
reg w13;    //: /sn:0 {0}(316,934)(140,934){1}
//: {2}(138,932)(138,816){3}
//: {4}(138,812)(138,761)(314,761){5}
//: {6}(136,814)(56,814){7}
//: {8}(138,936)(138,1433)(316,1433){9}
reg w94;    //: /sn:0 {0}(693,1376)(663,1376)(663,1431)(610,1431){1}
reg w5;    //: /sn:0 {0}(636,723)(703,723)(703,676)(718,676){1}
reg w48;    //: /sn:0 {0}(648,275)(683,275)(683,215)(822,215){1}
reg w47;    //: /sn:0 {0}(822,199)(667,199)(667,231)(648,231){1}
reg w107;    //: /sn:0 {0}(693,1312)(642,1312)(642,1271)(620,1271){1}
reg w145;    //: /sn:0 {0}(981,49)(1053,49)(1053,131)(1085,131){1}
reg w39;    //: /sn:0 {0}(309,404)(236,404){1}
//: {2}(234,402)(234,253){3}
//: {4}(236,251)(310,251){5}
//: {6}(234,249)(234,100){7}
//: {8}(236,98)(310,98){9}
//: {10}(232,98)(118,98)(118,175)(63,175){11}
//: {12}(234,406)(234,524){13}
//: {14}(236,526)(312,526){15}
//: {16}(234,528)(234,1543){17}
//: {18}(236,1545)(319,1545){19}
//: {20}(234,1547)(234,1698){21}
//: {22}(236,1700)(317,1700){23}
//: {24}(234,1702)(234,1897){25}
//: {26}(236,1899)(319,1899){27}
//: {28}(234,1901)(234,2051)(319,2051){29}
wire w32;    //: /sn:0 {0}(462,342)(462,388)(385,388){1}
wire w160;    //: /sn:0 {0}(1296,540)(1296,635)(1196,635){1}
wire w96;    //: /sn:0 {0}(459,1987)(459,2035)(402,2035){1}
wire w73;    //: /sn:0 {0}(954,1029)(873,1029)(873,1044)(842,1044){1}
wire w122;    //: /sn:0 {0}(1180,147)(1204,147){1}
//: {2}(1208,147)(1251,147)(1251,151)(1259,151){3}
//: {4}(1206,145)(1206,65){5}
wire [9:0] w141;    //: /sn:0 {0}(#:487,1722)(521,1722){1}
wire w56;    //: /sn:0 {0}(830,612)(871,612)(871,579){1}
wire w16;    //: /sn:0 {0}(485,469)(485,526)(388,526){1}
wire w179;    //: /sn:0 {0}(481,1707)(434,1707)(434,1700)(408,1700){1}
wire w81;    //: /sn:0 {0}(954,949)(923,949)(923,916)(842,916){1}
wire w19;    //: /sn:0 {0}(388,478)(410,478)(410,469){1}
wire w182;    //: /sn:0 {0}(408,1652)(456,1652)(456,1677)(481,1677){1}
wire w180;    //: /sn:0 {0}(481,1697)(439,1697)(439,1684)(408,1684){1}
wire w181;    //: /sn:0 {0}(481,1687)(447,1687)(447,1668)(408,1668){1}
wire w127;    //: /sn:0 {0}(1180,179)(1247,179){1}
wire w128;    //: /sn:0 {0}(393,990)(443,990)(443,956){1}
wire w104;    //: /sn:0 {0}(864,1263)(864,1280)(812,1280){1}
wire w75;    //: /sn:0 {0}(954,1009)(864,1009)(864,1012)(842,1012){1}
wire w67;    //: /sn:0 {0}(395,1883)(455,1883)(455,1835){1}
wire w54;    //: /sn:0 {0}(395,1497)(414,1497)(414,1481){1}
wire w119;    //: /sn:0 {0}(807,1537)(837,1537)(837,1525){1}
wire w176;    //: /sn:0 {0}(406,1321)(443,1321)(443,1285){1}
wire w174;    //: /sn:0 {0}(481,1727)(423,1727)(423,1732)(408,1732){1}
wire w124;    //: /sn:0 {0}(1247,212)(1193,212)(1193,211)(1180,211){1}
wire w20;    //: /sn:0 {0}(407,190)(407,203)(386,203){1}
wire w23;    //: /sn:0 {0}(486,190)(486,251)(386,251){1}
wire w82;    //: /sn:0 {0}(954,939)(932,939)(932,900)(842,900){1}
wire w158;    //: /sn:0 {0}(408,1780)(447,1780)(447,1757)(481,1757){1}
wire w125;    //: /sn:0 {0}(1247,196)(1192,196)(1192,195)(1180,195){1}
wire w74;    //: /sn:0 {0}(842,1028)(860,1028)(860,1019)(954,1019){1}
wire w8;    //: /sn:0 {0}(386,50)(409,50)(409,36){1}
wire w35;    //: /sn:0 {0}(385,436)(537,436)(537,343){1}
wire w103;    //: /sn:0 {0}(886,1263)(886,1296)(812,1296){1}
wire w163;    //: /sn:0 {0}(1196,587)(1239,587)(1239,539){1}
wire w71;    //: /sn:0 {0}(954,1049)(898,1049)(898,1076)(842,1076){1}
wire w101;    //: /sn:0 {0}(923,1263)(923,1328)(812,1328){1}
wire w22;    //: /sn:0 {0}(459,190)(459,235)(386,235){1}
wire w17;    //: /sn:0 {0}(458,469)(458,510)(388,510){1}
wire w53;    //: /sn:0 {0}(395,1513)(436,1513)(436,1481){1}
wire w117;    //: /sn:0 {0}(807,1569)(883,1569)(883,1525){1}
wire w113;    //: /sn:0 {0}(807,1633)(975,1633)(975,1525){1}
wire w83;    //: /sn:0 {0}(954,929)(941,929)(941,884)(842,884){1}
wire w77;    //: /sn:0 {0}(954,989)(881,989)(881,980)(842,980){1}
wire w115;    //: /sn:0 {0}(807,1601)(929,1601)(929,1525){1}
wire w78;    //: /sn:0 {0}(954,979)(891,979)(891,964)(842,964){1}
wire w10;    //: /sn:0 {0}(461,36)(461,82)(386,82){1}
wire w27;    //: /sn:0 {0}(390,633)(412,633)(412,612){1}
wire w95;    //: /sn:0 {0}(481,1987)(481,2051)(402,2051){1}
wire w52;    //: /sn:0 {0}(459,1482)(459,1529)(395,1529){1}
wire w178;    //: /sn:0 {0}(408,1716)(453,1716)(453,1717)(481,1717){1}
wire w80;    //: /sn:0 {0}(954,959)(912,959)(912,932)(842,932){1}
wire w29;    //: /sn:0 {0}(915,580)(915,644)(830,644){1}
wire w42;    //: /sn:0 {0}(886,135)(909,135)(909,118){1}
wire w175;    //: /sn:0 {0}(406,1337)(460,1337)(460,1285){1}
wire [15:0] w60;    //: /sn:0 {0}(989,1004)(#:960,1004){1}
wire w112;    //: /sn:0 {0}(807,1649)(998,1649)(998,1525){1}
wire w135;    //: /sn:0 {0}(393,1144)(443,1144)(443,1115){1}
wire w69;    //: /sn:0 {0}(395,1851)(414,1851)(414,1835){1}
wire w51;    //: /sn:0 {0}(481,1482)(481,1545)(395,1545){1}
wire w129;    //: /sn:0 {0}(392,838)(465,838)(465,790){1}
wire w97;    //: /sn:0 {0}(436,1987)(436,2019)(402,2019){1}
wire w114;    //: /sn:0 {0}(807,1617)(952,1617)(952,1525){1}
wire w177;    //: /sn:0 {0}(426,1285)(426,1305)(406,1305){1}
wire w66;    //: /sn:0 {0}(395,1899)(478,1899)(478,1836){1}
wire w64;    //: /sn:0 {0}(954,1079)(940,1079)(940,1124)(842,1124){1}
wire w34;    //: /sn:0 {0}(513,343)(513,420)(385,420){1}
wire w76;    //: /sn:0 {0}(954,999)(864,999)(864,996)(842,996){1}
wire w21;    //: /sn:0 {0}(386,219)(434,219)(434,190){1}
wire w102;    //: /sn:0 {0}(905,1263)(905,1312)(812,1312){1}
wire w157;    //: /sn:0 {0}(408,1796)(454,1796)(454,1767)(481,1767){1}
wire w31;    //: /sn:0 {0}(437,342)(437,372)(385,372){1}
wire w100;    //: /sn:0 {0}(812,1344)(947,1344)(947,1263){1}
wire w130;    //: /sn:0 {0}(392,822)(443,822)(443,790){1}
wire w161;    //: /sn:0 {0}(1196,619)(1276,619)(1276,541){1}
wire w132;    //: /sn:0 {0}(393,974)(417,974)(417,956){1}
wire w140;    //: /sn:0 {0}(1180,115)(1235,115){1}
//: {2}(1239,115)(1248,115)(1248,131)(1259,131){3}
//: {4}(1237,113)(1237,64){5}
wire w25;    //: /sn:0 {0}(390,665)(464,665)(464,612){1}
wire w116;    //: /sn:0 {0}(807,1585)(906,1585)(906,1525){1}
wire w98;    //: /sn:0 {0}(418,1987)(418,2003)(402,2003){1}
wire w65;    //: /sn:0 {0}(954,1069)(925,1069)(925,1108)(842,1108){1}
wire w118;    //: /sn:0 {0}(807,1553)(860,1553)(860,1525){1}
wire w18;    //: /sn:0 {0}(434,469)(434,494)(388,494){1}
wire w164;    //: /sn:0 {0}(1196,571)(1222,571)(1222,539){1}
wire w162;    //: /sn:0 {0}(1196,603)(1257,603)(1257,540){1}
wire w30;    //: /sn:0 {0}(410,342)(410,356)(385,356){1}
wire w68;    //: /sn:0 {0}(395,1867)(432,1867)(432,1835){1}
wire w123;    //: /sn:0 {0}(1180,131)(1218,131){1}
//: {2}(1222,131)(1237,131)(1237,141)(1259,141){3}
//: {4}(1220,129)(1220,119)(1221,119)(1221,65){5}
wire w165;    //: /sn:0 {0}(408,1764)(437,1764)(437,1747)(481,1747){1}
wire w137;    //: /sn:0 {0}(1247,228)(1194,228)(1194,227)(1180,227){1}
wire w11;    //: /sn:0 {0}(488,36)(488,98)(386,98){1}
wire w57;    //: /sn:0 {0}(830,596)(850,596)(850,580){1}
wire w136;    //: /sn:0 {0}(393,1128)(417,1128)(417,1115){1}
wire w139;    //: /sn:0 {0}(1180,163)(1187,163){1}
//: {2}(1191,163)(1245,163)(1245,161)(1259,161){3}
//: {4}(1189,161)(1189,65){5}
wire w173;    //: /sn:0 {0}(408,1748)(428,1748)(428,1737)(481,1737){1}
wire w70;    //: /sn:0 {0}(954,1059)(913,1059)(913,1092)(842,1092){1}
wire w72;    //: /sn:0 {0}(954,1039)(886,1039)(886,1060)(842,1060){1}
wire w33;    //: /sn:0 {0}(489,342)(489,404)(385,404){1}
wire w131;    //: /sn:0 {0}(392,806)(422,806)(422,790){1}
wire [3:0] w143;    //: /sn:0 {0}(#:1265,146)(1317,146){1}
wire w9;    //: /sn:0 {0}(436,36)(436,66)(386,66){1}
wire w79;    //: /sn:0 {0}(954,969)(902,969)(902,948)(842,948){1}
wire w55;    //: /sn:0 {0}(893,579)(893,628)(830,628){1}
wire w26;    //: /sn:0 {0}(440,612)(440,649)(390,649){1}
//: enddecls

  //: joint g165 (w0) @(221, 1006) /w:[ 22 21 -1 24 ]
  //: joint g8 (w0) @(221, 267) /w:[ 12 14 -1 11 ]
  //: SWITCH g140 (w120) @(717,1705) /sn:0 /w:[ 0 ] /st:0 /dn:0
  //: LED g37 (w34) @(513,336) /sn:0 /w:[ 0 ] /type:0
  //: joint g13 (w38) @(250, 82) /w:[ 28 -1 30 27 ]
  //: joint g55 (w36) @(280, 633) /w:[ 4 6 -1 3 ]
  //: LED g139 (w112) @(998,1518) /sn:0 /w:[ 1 ] /type:0
  //: joint g111 (w1) @(209, 1931) /w:[ 38 37 -1 40 ]
  //: LED g218 (w160) @(1296,533) /sn:0 /w:[ 0 ] /type:0
  //: joint g176 (w7) @(166, 1038) /w:[ 10 9 -1 12 ]
  H7402 g1 (.B4(w3), .B3(w2), .B2(w1), .B1(w0), .A4(w39), .A3(w38), .A2(w37), .A1(w36), .Y4(w23), .Y3(w22), .Y2(w21), .Y1(w20));   //: @(311, 187) /sz:(74, 144) /sn:0 /p:[ Li0>0 Li1>17 Li2>13 Li3>13 Li4>5 Li5>25 Li6>17 Li7>17 Ro0<1 Ro1<1 Ro2<0 Ro3<1 ]
  //: SWITCH D1 (w133) @(34,976) /w:[ 0 ] /st:0 /dn:0
  //: SWITCH A (w43) @(632,44) /w:[ 0 ] /st:1 /dn:0
  //: joint g11 (w36) @(280, 50) /w:[ 20 -1 22 19 ]
  //: SWITCH g130 (w99) @(593,1466) /sn:0 /w:[ 1 ] /st:0 /dn:0
  //: SWITCH C3 (w13) @(39,814) /w:[ 7 ] /st:0 /dn:0
  //: LED g50 (w26) @(440,605) /sn:0 /w:[ 0 ] /type:0
  //: joint g223 (w0) @(221, 1353) /w:[ 30 29 -1 32 ]
  //: LED g197 (w127) @(1254,179) /sn:0 /R:3 /w:[ 1 ] /type:0
  //: LED g132 (w119) @(837,1518) /sn:0 /w:[ 1 ] /type:0
  //: joint g113 (w3) @(180, 1963) /w:[ 18 17 -1 20 ]
  //: SWITCH A6 (w40) @(49,460) /w:[ 0 ] /st:0 /dn:0
  //: joint g19 (w36) @(280, 203) /w:[ 16 18 -1 15 ]
  //: LED g150 (w129) @(465,783) /sn:0 /w:[ 1 ] /type:0
  //: SWITCH g146 (w110) @(604,1688) /sn:0 /w:[ 0 ] /st:0 /dn:0
  //: SWITCH A2 (w37) @(46,91) /w:[ 23 ] /st:1 /dn:0
  //: SWITCH g115 (w59) @(131,2162) /sn:0 /w:[ 0 ] /st:0 /dn:0
  //: LED g38 (w35) @(537,336) /sn:0 /w:[ 1 ] /type:0
  //: LED g75 (w56) @(871,572) /sn:0 /w:[ 1 ] /type:0
  //: joint g227 (w12) @(152, 1208) /w:[ 14 13 -1 16 ]
  H7421 g169 (.A1(w36), .A2(w37), .B1(w0), .B2(w1), .C1(w7), .C2(w12), .D1(w133), .D2(w134), .Y1(w136), .Y2(w135));   //: @(318, 1112) /sz:(74, 144) /sn:0 /p:[ Li0>31 Li1>31 Li2>27 Li3>27 Li4>15 Li5>15 Li6>5 Li7>5 Ro0<0 Ro1<0 ]
  H7420 g160 (.A1(w36), .A2(w37), .B1(w0), .B2(w1), .C1(w7), .C2(w12), .D1(w133), .D2(w134), .Y1(w132), .Y2(w128));   //: @(318, 958) /sz:(74, 144) /sn:0 /p:[ Li0>27 Li1>27 Li2>23 Li3>23 Li4>11 Li5>11 Li6>3 Li7>3 Ro0<0 Ro1<0 ]
  //: LED g135 (w116) @(906,1518) /sn:0 /w:[ 1 ] /type:0
  //: LED g31 (w20) @(407,183) /sn:0 /w:[ 0 ] /type:0
  //: joint g20 (w37) @(266, 219) /w:[ 16 18 -1 15 ]
  //: SWITCH g124 (w107) @(603,1271) /sn:0 /w:[ 1 ] /st:0 /dn:0
  //: LED g230 (w176) @(443,1278) /sn:0 /w:[ 1 ] /type:0
  //: LED g39 (w18) @(434,462) /sn:0 /w:[ 0 ] /type:0
  //: SWITCH g68 (w58) @(618,543) /sn:0 /w:[ 0 ] /st:0 /dn:0
  //: SWITCH g195 (w154) @(963,359) /sn:0 /w:[ 0 ] /st:1 /dn:0
  //: LED g205 (w122) @(1206,58) /sn:0 /w:[ 5 ] /type:0
  //: joint g179 (w134) @(77, 1086) /w:[ 2 1 -1 4 ]
  H7430 g52 (.A(w43), .B(w44), .C(w45), .D(w46), .E(w47), .F(w48), .G(w49), .H(w50), .Y(w42));   //: @(823, 119) /sz:(62, 144) /sn:0 /p:[ Li0>1 Li1>0 Li2>0 Li3>0 Li4>0 Li5>1 Li6>1 Li7>1 Ro0<0 ]
  //: joint g107 (w37) @(266, 1867) /w:[ 46 45 -1 48 ]
  //: LED g231 (w175) @(460,1278) /sn:0 /w:[ 1 ] /type:0
  //: joint g221 (w37) @(266, 1321) /w:[ 34 33 -1 36 ]
  //: LED g201 (w140) @(1237,57) /sn:0 /w:[ 5 ] /type:0
  //: joint g14 (w39) @(234, 98) /w:[ 8 -1 10 7 ]
  //: joint g47 (w1) @(209, 558) /w:[ 8 10 -1 7 ]
  //: joint g44 (w37) @(266, 494) /w:[ 8 10 -1 7 ]
  //: SWITCH C (w45) @(630,135) /w:[ 1 ] /st:1 /dn:0
  //: joint g84 (w0) @(221, 1561) /w:[ 34 33 -1 36 ]
  //: LED g105 (w95) @(481,1980) /sn:0 /w:[ 0 ] /type:0
  //: LED g236 (w141) @(528,1722) /sn:0 /R:3 /w:[ 1 ] /type:1
  //: joint g23 (w3) @(181, 315) /w:[ 1 2 -1 8 ]
  H74163 g116 (.A(w105), .B(w106), .C(w107), .D(w108), ._CLR(w92), .ENP(w93), .ENT(w94), ._LOAD(w99), .CLK(w91), .QA(w104), .QB(w103), .QC(w102), .QD(w101), .RCO(w100));   //: @(694, 1264) /sz:(117, 160) /sn:0 /p:[ Li0>0 Li1>0 Li2>0 Li3>1 Li4>0 Li5>0 Li6>0 Li7>0 Bi0>1 Ro0<1 Ro1<1 Ro2<1 Ro3<1 Ro4<0 ]
  //: LED g40 (w17) @(458,462) /sn:0 /w:[ 0 ] /type:0
  //: SWITCH A1 (w36) @(46,50) /w:[ 23 ] /st:0 /dn:0
  H7432 g54 (.A1(w36), .A2(w37), .A3(w38), .A4(w39), .B1(w0), .B2(w1), .B3(w2), .B4(w3), .Y1(w54), .Y2(w53), .Y3(w52), .Y4(w51));   //: @(320, 1481) /sz:(74, 144) /sn:0 /p:[ Li0>39 Li1>39 Li2>0 Li3>19 Li4>35 Li5>35 Li6>27 Li7>15 Ro0<0 Ro1<0 Ro2<1 Ro3<1 ]
  //: SWITCH g93 (w84) @(620,867) /sn:0 /w:[ 0 ] /st:0 /dn:0
  //: joint g167 (w7) @(166, 902) /w:[ 1 2 -1 8 ]
  //: joint g46 (w0) @(221, 542) /w:[ 8 10 -1 7 ]
  //: LED g26 (w9) @(436,29) /sn:0 /w:[ 0 ] /type:0
  H7400 g0 (.B4(w3), .B3(w2), .B2(w1), .B1(w0), .A4(w39), .A3(w38), .A2(w37), .A1(w36), .Y4(w11), .Y3(w10), .Y2(w9), .Y1(w8));   //: @(311, 34) /sz:(74, 144) /sn:0 /p:[ Li0>5 Li1>21 Li2>17 Li3>17 Li4>9 Li5>29 Li6>21 Li7>21 Ro0<1 Ro1<1 Ro2<1 Ro3<0 ]
  //: joint g228 (w13) @(138, 934) /w:[ 1 2 -1 8 ]
  //: joint g224 (w1) @(209, 1368) /w:[ 30 29 -1 32 ]
  //: LED g136 (w115) @(929,1518) /sn:0 /w:[ 1 ] /type:0
  //: joint g233 (w36) @(280, 1652) /w:[ 42 41 -1 44 ]
  //: SWITCH g190 (w151) @(964,186) /sn:0 /w:[ 1 ] /st:0 /dn:0
  //: joint g173 (w37) @(266, 1143) /w:[ 30 29 -1 32 ]
  //: SWITCH _G2 (w167) @(991,578) /w:[ 0 ] /st:0 /dn:0
  //: joint g61 (w2) @(195, 713) /w:[ 8 10 -1 7 ]
  //: joint g220 (w36) @(280, 1305) /w:[ 34 33 -1 36 ]
  //: joint g3 (w36) @(280, 356) /w:[ 12 14 -1 11 ]
  //: LED g34 (w30) @(410,335) /sn:0 /w:[ 0 ] /type:0
  //: joint g86 (w2) @(195, 1593) /w:[ 26 25 -1 28 ]
  //: joint g110 (w0) @(221, 1915) /w:[ 38 37 -1 40 ]
  //: LED g65 (w52) @(459,1475) /sn:0 /w:[ 0 ] /type:0
  //: joint g59 (w0) @(221, 681) /w:[ 4 6 -1 3 ]
  //: SWITCH F (w48) @(631,275) /w:[ 0 ] /st:1 /dn:0
  H7411 g147 (.A1(w36), .A2(w37), .A3(w38), .B1(w0), .B2(w1), .B3(w2), .C1(w7), .C2(w12), .C3(w13), .Y1(w131), .Y2(w130), .Y3(w129));   //: @(317, 790) /sz:(74, 160) /sn:0 /p:[ Li0>0 Li1>0 Li2>9 Li3>0 Li4>0 Li5>5 Li6>0 Li7>0 Li8>0 Ro0<0 Ro1<0 Ro2<0 ]
  //: joint g156 (w2) @(195, 887) /w:[ 4 6 -1 3 ]
  //: joint g153 (w38) @(250, 838) /w:[ 8 10 -1 7 ]
  //: SWITCH g98 (w89) @(620,1049) /sn:0 /w:[ 0 ] /st:0 /dn:0
  //: joint g16 (w1) @(209, 130) /w:[ 16 -1 18 15 ]
  //: SWITCH g96 (w87) @(620,977) /sn:0 /w:[ 0 ] /st:0 /dn:0
  //: SWITCH g183 (w144) @(964,18) /sn:0 /w:[ 0 ] /st:0 /dn:0
  //: SWITCH g122 (w105) @(602,1212) /sn:0 /w:[ 1 ] /st:0 /dn:0
  //: SWITCH g78 (w4) @(704,768) /sn:0 /w:[ 1 ] /st:0 /dn:0
  //: joint g87 (w3) @(181, 1609) /w:[ 14 13 -1 16 ]
  //: SWITCH g129 (w94) @(593,1431) /sn:0 /w:[ 1 ] /st:0 /dn:0
  //: LED g171 (w135) @(443,1108) /sn:0 /w:[ 1 ] /type:0
  //: SWITCH g69 (w24) @(617,574) /sn:0 /w:[ 0 ] /st:0 /dn:0
  //: SWITCH g143 (w109) @(604,1593) /sn:0 /w:[ 0 ] /st:0 /dn:0
  //: LED g119 (w102) @(905,1256) /sn:0 /w:[ 0 ] /type:0
  //: joint g15 (w0) @(221, 114) /w:[ 16 -1 18 15 ]
  //: SWITCH C2 (w12) @(38,772) /w:[ 7 ] /st:0 /dn:0
  //: LED g162 (w128) @(443,949) /sn:0 /w:[ 1 ] /type:0
  H74175 g131 (.D1(w111), .D2(w121), .D3(w109), .D4(w90), ._PRE(w63), ._CLR(w110), .CLK(w120), .Q1(w119), .Q2(w118), .Q3(w117), .Q4(w116), ._Q1(w115), ._Q2(w114), ._Q3(w113), ._Q4(w112));   //: @(701, 1521) /sz:(105, 144) /sn:0 /p:[ Li0>1 Li1>0 Li2>1 Li3>1 Li4>1 Li5>1 Bi0>1 Ro0<0 Ro1<0 Ro2<0 Ro3<0 Ro4<0 Ro5<0 Ro6<0 Ro7<0 ]
  //: SWITCH g127 (w92) @(593,1366) /sn:0 /w:[ 1 ] /st:1 /dn:0
  H7474 g67 (.D1(w58), ._PRE1(w24), ._CLR1(w15), .D2(w14), ._PRE2(w6), ._CLR2(w5), .CLK(w4), .Q1(w57), ._Q1(w56), .Q2(w55), ._Q2(w29));   //: @(719, 580) /sz:(110, 124) /sn:0 /p:[ Li0>1 Li1>1 Li2>1 Li3>1 Li4>1 Li5>1 Bi0>0 Ro0<0 Ro1<0 Ro2<1 Ro3<1 ]
  //: joint g43 (w36) @(280, 478) /w:[ 8 10 -1 7 ]
  //: joint g62 (w3) @(181, 590) /w:[ 10 9 -1 12 ]
  //: LED g88 (w69) @(414,1828) /sn:0 /w:[ 1 ] /type:0
  //: LED g104 (w96) @(459,1980) /sn:0 /w:[ 0 ] /type:0
  //: SWITCH g188 (w149) @(964,155) /sn:0 /w:[ 0 ] /st:0 /dn:0
  //: LED g63 (w54) @(414,1474) /sn:0 /w:[ 1 ] /type:0
  //: LED g138 (w113) @(975,1518) /sn:0 /w:[ 1 ] /type:0
  //: SWITCH Cn (w126) @(990,841) /w:[ 0 ] /st:0 /dn:0
  //: joint g109 (w39) @(234, 1899) /w:[ 26 25 -1 28 ]
  //: joint g175 (w1) @(209, 1175) /w:[ 26 25 -1 28 ]
  //: joint g234 (w37) @(266, 1668) /w:[ 42 41 -1 44 ]
  //: LED g133 (w118) @(860,1518) /sn:0 /w:[ 1 ] /type:0
  //: joint g5 (w37) @(266, 372) /w:[ 12 14 -1 11 ]
  //: joint g56 (w37) @(266, 649) /w:[ 4 6 -1 3 ]
  //: SWITCH g95 (w86) @(620,941) /sn:0 /w:[ 0 ] /st:0 /dn:0
  //: LED g24 (w19) @(410,462) /sn:0 /w:[ 1 ] /type:0
  //: joint g85 (w1) @(209, 1577) /w:[ 34 33 -1 36 ]
  H74154 g92 (.A(w84), .B(w85), .C(w86), .D(w87), ._G1(w88), ._G2(w89), ._Y1(w83), ._Y2(w82), ._Y3(w81), ._Y4(w80), ._Y5(w79), ._Y6(w78), ._Y7(w77), ._Y8(w76), ._Y9(w75), ._Y10(w74), ._Y11(w73), ._Y12(w72), ._Y13(w71), ._Y14(w70), ._Y15(w65), ._Y16(w64));   //: @(736, 868) /sz:(105, 272) /sn:0 /p:[ Li0>1 Li1>0 Li2>1 Li3>1 Li4>1 Li5>1 Ro0<1 Ro1<1 Ro2<1 Ro3<1 Ro4<1 Ro5<1 Ro6<1 Ro7<1 Ro8<1 Ro9<0 Ro10<1 Ro11<1 Ro12<1 Ro13<1 Ro14<1 Ro15<1 ]
  //: LED g214 (w164) @(1222,532) /sn:0 /w:[ 1 ] /type:0
  //: SWITCH g210 (w169) @(991,756) /w:[ 0 ] /st:0 /dn:0
  //: joint g60 (w1) @(209, 697) /w:[ 4 6 -1 3 ]
  H74157 g101 (.A1(w36), .A2(w37), .A3(w38), .A4(w39), .B1(w0), .B2(w1), .B3(w2), .B4(w3), ._G(w61), .S(w59), .Y1(w98), .Y2(w97), .Y3(w96), .Y4(w95));   //: @(320, 1987) /sz:(81, 176) /sn:0 /p:[ Li0>49 Li1>49 Li2>41 Li3>29 Li4>41 Li5>41 Li6>33 Li7>21 Li8>0 Li9>1 Ro0<1 Ro1<1 Ro2<1 Ro3<1 ]
  //: SWITCH g185 (w146) @(964,81) /sn:0 /w:[ 0 ] /st:0 /dn:0
  //: SWITCH g126 (w91) @(712,1495) /sn:0 /w:[ 0 ] /st:0 /dn:0
  //: LED g35 (w33) @(489,335) /sn:0 /w:[ 0 ] /type:0
  //: LED g170 (w136) @(417,1108) /sn:0 /w:[ 1 ] /type:0
  //: joint g204 (w123) @(1220, 131) /w:[ 2 4 1 -1 ]
  //: SWITCH C1 (w7) @(39,729) /w:[ 7 ] /st:1 /dn:0
  //: joint g235 (w38) @(250, 1684) /w:[ 34 33 -1 36 ]
  //: SWITCH E (w47) @(631,231) /w:[ 1 ] /st:1 /dn:0
  //: SWITCH B3 (w2) @(46,313) /w:[ 23 ] /st:0 /dn:0
  //: LED g66 (w51) @(481,1475) /sn:0 /w:[ 0 ] /type:0
  //: SWITCH g97 (w88) @(620,1013) /sn:0 /w:[ 0 ] /st:0 /dn:0
  //: LED g120 (w101) @(923,1256) /sn:0 /w:[ 0 ] /type:0
  //: SWITCH g184 (w145) @(964,49) /sn:0 /w:[ 0 ] /st:0 /dn:0
  //: joint g18 (w3) @(181, 162) /w:[ 4 -1 6 3 ]
  //: joint g12 (w37) @(266, 66) /w:[ 20 -1 22 19 ]
  //: joint g226 (w7) @(166, 1192) /w:[ 14 13 -1 16 ]
  H7427 g219 (.A1(w36), .A2(w37), .A3(w38), .B1(w0), .B2(w1), .B3(w2), .C1(w7), .C2(w12), .C3(w13), .Y1(w177), .Y2(w176), .Y3(w175));   //: @(317, 1289) /sz:(88, 160) /sn:0 /p:[ Li0>35 Li1>35 Li2>5 Li3>31 Li4>31 Li5>0 Li6>17 Li7>17 Li8>9 Ro0<1 Ro1<0 Ro2<0 ]
  //: joint g108 (w38) @(250, 1883) /w:[ 38 37 -1 40 ]
  //: SWITCH A4 (w39) @(46,175) /w:[ 11 ] /st:1 /dn:0
  //: SWITCH g191 (w28) @(964,296) /sn:0 /w:[ 0 ] /st:1 /dn:0
  //: SWITCH _G1 (w159) @(991,536) /w:[ 1 ] /st:0 /dn:0
  //: LED g134 (w117) @(883,1518) /sn:0 /w:[ 1 ] /type:0
  assign w141 = {w157, w158, w165, w173, w174, w178, w179, w180, w181, w182}; //: CONCAT g237  @(486,1722) /sn:0 /w:[ 0 1 1 1 1 0 1 0 0 0 1 ] /dr:1 /tp:1 /drp:1
  H7408 g4 (.A1(w36), .A2(w37), .A3(w38), .A4(w39), .B1(w0), .B2(w1), .B3(w2), .B4(w3), .Y1(w19), .Y2(w18), .Y3(w17), .Y4(w16));   //: @(313, 462) /sz:(74, 144) /sn:0 /p:[ Li0>9 Li1>9 Li2>17 Li3>15 Li4>9 Li5>9 Li6>13 Li7>11 Ro0<0 Ro1<1 Ro2<1 Ro3<1 ]
  //: joint g154 (w0) @(221, 854) /w:[ 1 2 -1 20 ]
  //: joint g58 (w39) @(234, 526) /w:[ 14 13 -1 16 ]
  //: SWITCH g186 (w147) @(964,114) /sn:0 /w:[ 0 ] /st:0 /dn:0
  //: joint g112 (w2) @(195, 1947) /w:[ 30 29 -1 32 ]
  //: LED g76 (w55) @(893,572) /sn:0 /w:[ 0 ] /type:0
  //: SWITCH g211 (w170) @(991,797) /w:[ 1 ] /st:0 /dn:0
  //: joint g157 (w7) @(166, 729) /w:[ 4 -1 6 3 ]
  //: joint g238 (w39) @(234, 1700) /w:[ 22 21 -1 24 ]
  //: SWITCH A3 (w38) @(46,134) /w:[ 31 ] /st:0 /dn:0
  //: joint g163 (w36) @(280, 974) /w:[ 26 25 -1 28 ]
  //: LED g64 (w53) @(436,1474) /sn:0 /w:[ 1 ] /type:0
  //: SWITCH D2 (w134) @(34,1021) /w:[ 0 ] /st:0 /dn:0
  //: joint g166 (w1) @(209, 1022) /w:[ 22 21 -1 24 ]
  //: LED g121 (w100) @(947,1256) /sn:0 /w:[ 1 ] /type:0
  //: joint g206 (w122) @(1206, 147) /w:[ 2 4 1 -1 ]
  //: LED g28 (w11) @(488,29) /sn:0 /w:[ 0 ] /type:0
  //: SWITCH G (w49) @(631,322) /w:[ 0 ] /st:1 /dn:0
  //: joint g225 (w2) @(195, 1385) /w:[ 1 2 -1 24 ]
  //: SWITCH B2 (w1) @(46,272) /w:[ 19 ] /st:0 /dn:0
  //: joint g6 (w38) @(250, 388) /w:[ 20 22 -1 19 ]
  //: joint g177 (w12) @(152, 1054) /w:[ 10 9 -1 12 ]
  //: SWITCH g192 (w62) @(964,324) /sn:0 /w:[ 0 ] /st:0 /dn:0
  //: joint g208 (w139) @(1189, 163) /w:[ 2 4 1 -1 ]
  //: joint g7 (w39) @(234, 404) /w:[ 1 2 -1 12 ]
  //: LED g53 (w42) @(909,111) /sn:0 /w:[ 1 ] /type:0
  //: LED g149 (w130) @(443,783) /sn:0 /w:[ 1 ] /type:0
  //: SWITCH B1 (w0) @(46,231) /w:[ 19 ] /st:0 /dn:0
  //: LED g207 (w139) @(1189,58) /sn:0 /w:[ 5 ] /type:0
  //: joint g48 (w2) @(195, 574) /w:[ 12 14 -1 11 ]
  //: LED g200 (w137) @(1254,228) /sn:0 /R:3 /w:[ 0 ] /type:0
  //: joint g17 (w2) @(195, 146) /w:[ 20 -1 22 19 ]
  //: LED g25 (w8) @(409,29) /sn:0 /w:[ 1 ] /type:0
  //: LED g29 (w23) @(486,183) /sn:0 /w:[ 0 ] /type:0
  //: joint g106 (w36) @(280, 1851) /w:[ 46 45 -1 48 ]
  //: joint g83 (w39) @(234, 1545) /w:[ 18 17 -1 20 ]
  //: joint g174 (w0) @(221, 1159) /w:[ 26 25 -1 28 ]
  //: LED g100 (w60) @(996,1004) /sn:0 /R:3 /w:[ 0 ] /type:1
  //: SWITCH g94 (w85) @(620,905) /sn:0 /w:[ 1 ] /st:0 /dn:0
  //: joint g80 (w36) @(280, 1497) /w:[ 38 37 -1 40 ]
  //: SWITCH g193 (w152) @(963,422) /sn:0 /w:[ 1 ] /st:0 /dn:0
  //: joint g202 (w140) @(1237, 115) /w:[ 2 4 1 -1 ]
  H7442 g232 (.A3(w39), .A2(w38), .A1(w37), .A0(w36), ._Y9(w157), ._Y8(w158), ._Y7(w165), ._Y6(w173), ._Y5(w174), ._Y4(w178), ._Y3(w179), ._Y2(w180), ._Y1(w181), ._Y0(w182));   //: @(318, 1636) /sz:(89, 175) /sn:0 /p:[ Li0>23 Li1>35 Li2>43 Li3>43 Ro0<0 Ro1<0 Ro2<0 Ro3<0 Ro4<1 Ro5<0 Ro6<1 Ro7<1 Ro8<1 Ro9<0 ]
  //: joint g21 (w38) @(250, 235) /w:[ 24 26 -1 23 ]
  //: SWITCH D (w46) @(631,183) /w:[ 1 ] /st:1 /dn:0
  //: joint g159 (w13) @(138, 814) /w:[ -1 4 6 3 ]
  //: joint g172 (w36) @(280, 1128) /w:[ 30 29 -1 32 ]
  //: LED g41 (w16) @(485,462) /sn:0 /w:[ 0 ] /type:0
  //: SWITCH g141 (w111) @(604,1537) /sn:0 /w:[ 0 ] /st:0 /dn:0
  //: joint g155 (w1) @(209, 870) /w:[ 1 2 -1 20 ]
  //: SWITCH g123 (w106) @(602,1241) /sn:0 /w:[ 1 ] /st:0 /dn:0
  //: joint g151 (w36) @(280, 806) /w:[ 1 2 -1 24 ]
  //: LED g90 (w67) @(455,1828) /sn:0 /w:[ 1 ] /type:0
  //: joint g222 (w38) @(250, 1337) /w:[ 4 6 -1 3 ]
  //: joint g82 (w38) @(250, 1529) /w:[ 1 2 -1 32 ]
  //: SWITCH B4 (w3) @(46,354) /w:[ 7 ] /st:0 /dn:0
  //: SWITCH g128 (w93) @(593,1399) /sn:0 /w:[ 1 ] /st:0 /dn:0
  //: LED g91 (w66) @(478,1829) /sn:0 /w:[ 1 ] /type:0
  //: LED g33 (w31) @(437,335) /sn:0 /w:[ 0 ] /type:0
  //: LED g49 (w27) @(412,605) /sn:0 /w:[ 1 ] /type:0
  //: LED g137 (w114) @(952,1518) /sn:0 /w:[ 1 ] /type:0
  //: LED g198 (w125) @(1254,196) /sn:0 /R:3 /w:[ 0 ] /type:0
  //: LED g51 (w25) @(464,605) /sn:0 /w:[ 1 ] /type:0
  //: SWITCH B (w44) @(631,91) /w:[ 1 ] /st:1 /dn:0
  //: joint g158 (w12) @(152, 745) /w:[ 4 -1 6 3 ]
  //: LED g89 (w68) @(432,1828) /sn:0 /w:[ 1 ] /type:0
  //: SWITCH A5 (w41) @(49,420) /w:[ 0 ] /st:0 /dn:0
  //: SWITCH _G3 (w168) @(991,619) /w:[ 1 ] /st:0 /dn:0
  //: LED g217 (w161) @(1276,534) /sn:0 /w:[ 1 ] /type:0
  H7404 g2 (.A6(w40), .A5(w41), .A4(w39), .A3(w38), .A2(w37), .A1(w36), .Y6(w35), .Y5(w34), .Y4(w33), .Y3(w32), .Y2(w31), .Y1(w30));   //: @(310, 340) /sz:(74, 112) /sn:0 /p:[ Li0>1 Li1>1 Li2>0 Li3>21 Li4>13 Li5>13 Ro0<0 Ro1<1 Ro2<1 Ro3<1 Ro4<1 Ro5<1 ]
  //: LED g77 (w29) @(915,573) /sn:0 /w:[ 0 ] /type:0
  //: LED g148 (w131) @(422,783) /sn:0 /w:[ 1 ] /type:0
  //: SWITCH g213 (w172) @(991,714) /w:[ 0 ] /st:0 /dn:0
  //: LED g203 (w123) @(1221,58) /sn:0 /w:[ 5 ] /type:0
  //: SWITCH g72 (w6) @(618,690) /sn:0 /w:[ 0 ] /st:0 /dn:0
  assign w60 = {w64, w65, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83}; //: CONCAT g99  @(959,1004) /sn:0 /w:[ 1 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 ] /dr:1 /tp:0 /drp:1
  //: LED g161 (w132) @(417,949) /sn:0 /w:[ 1 ] /type:0
  assign w143 = {w139, w122, w123, w140}; //: CONCAT g182  @(1264,146) /sn:0 /w:[ 0 3 3 3 3 ] /dr:1 /tp:0 /drp:1
  //: SWITCH g196 (w155) @(963,390) /sn:0 /w:[ 1 ] /st:0 /dn:0
  //: joint g152 (w37) @(266, 822) /w:[ 1 2 -1 24 ]
  //: LED g103 (w98) @(418,1980) /sn:0 /w:[ 0 ] /type:0
  //: SWITCH g189 (w150) @(964,218) /sn:0 /w:[ 1 ] /st:0 /dn:0
  //: joint g10 (w2) @(195, 299) /w:[ 16 18 -1 15 ]
  //: SWITCH g212 (w171) @(991,673) /w:[ 0 ] /st:0 /dn:0
  //: LED g199 (w124) @(1254,212) /sn:0 /R:3 /w:[ 0 ] /type:0
  //: LED g32 (w21) @(434,183) /sn:0 /w:[ 1 ] /type:0
  //: LED g27 (w10) @(461,29) /sn:0 /w:[ 0 ] /type:0
  //: SWITCH _G0 (w166) @(991,495) /w:[ 0 ] /st:0 /dn:0
  //: LED g102 (w97) @(436,1980) /sn:0 /w:[ 0 ] /type:0
  //: SWITCH g187 (w148) @(964,251) /sn:0 /w:[ 0 ] /st:0 /dn:0
  //: joint g9 (w1) @(209, 283) /w:[ 12 14 -1 11 ]
  //: joint g57 (w38) @(250, 665) /w:[ 12 14 -1 11 ]
  //: SWITCH g71 (w14) @(617,658) /sn:0 /w:[ 0 ] /st:0 /dn:0
  //: SWITCH g142 (w121) @(604,1565) /sn:0 /w:[ 1 ] /st:0 /dn:0
  //: SWITCH g73 (w5) @(619,723) /sn:0 /w:[ 0 ] /st:0 /dn:0
  //: SWITCH g145 (w63) @(604,1663) /sn:0 /w:[ 0 ] /st:0 /dn:0
  H7410 g42 (.A1(w36), .A2(w37), .A3(w38), .B1(w0), .B2(w1), .B3(w2), .C1(w7), .C2(w12), .C3(w13), .Y1(w27), .Y2(w26), .Y3(w25));   //: @(315, 617) /sz:(74, 160) /sn:0 /p:[ Li0>5 Li1>5 Li2>13 Li3>5 Li4>5 Li5>9 Li6>5 Li7>5 Li8>5 Ro0<0 Ro1<1 Ro2<0 ]
  H74181 g180 (._A0(w144), ._A1(w145), ._A2(w146), ._A3(w147), ._B0(w149), ._B1(w151), ._B2(w150), ._B3(w148), .Cn(w28), .M(w62), .S0(w154), .S1(w155), .S2(w152), .S3(w153), ._F0(w140), ._F1(w123), ._F2(w122), ._F3(w139), .AEB(w127), .CnP4(w125), ._G(w124), ._P(w137));   //: @(1086, 99) /sz:(93, 240) /sn:0 /p:[ Li0>1 Li1>1 Li2>1 Li3>1 Li4>1 Li5>0 Li6>0 Li7>1 Li8>1 Li9>1 Li10>1 Li11>0 Li12>0 Li13>1 Ro0<0 Ro1<0 Ro2<0 Ro3<0 Ro4<0 Ro5<1 Ro6<1 Ro7<1 ]
  //: LED g74 (w57) @(850,573) /sn:0 /w:[ 1 ] /type:0
  //: joint g168 (w12) @(152, 918) /w:[ 1 2 -1 8 ]
  //: LED g181 (w143) @(1324,146) /sn:0 /R:3 /w:[ 1 ] /type:2
  H7486 g79 (.A1(w36), .A2(w37), .A3(w38), .A4(w39), .B1(w0), .B2(w1), .B3(w2), .B4(w3), .Y1(w69), .Y2(w68), .Y3(w67), .Y4(w66));   //: @(320, 1835) /sz:(74, 144) /sn:0 /p:[ Li0>47 Li1>47 Li2>39 Li3>27 Li4>39 Li5>39 Li6>31 Li7>19 Ro0<0 Ro1<0 Ro2<0 Ro3<0 ]
  //: SWITCH H (w50) @(631,368) /w:[ 0 ] /st:1 /dn:0
  //: LED g117 (w104) @(864,1256) /sn:0 /w:[ 0 ] /type:0
  //: SWITCH g194 (w153) @(963,455) /sn:0 /w:[ 0 ] /st:1 /dn:0
  //: LED g215 (w163) @(1239,532) /sn:0 /w:[ 1 ] /type:0
  //: LED g36 (w32) @(462,335) /sn:0 /w:[ 0 ] /type:0
  //: LED g216 (w162) @(1257,533) /sn:0 /w:[ 1 ] /type:0
  //: joint g178 (w133) @(91, 1070) /w:[ 2 1 -1 4 ]
  //: SWITCH g144 (w90) @(604,1622) /sn:0 /w:[ 0 ] /st:0 /dn:0
  //: SWITCH g125 (w108) @(602,1300) /sn:0 /w:[ 0 ] /st:0 /dn:0
  //: joint g81 (w37) @(266, 1513) /w:[ 38 37 -1 40 ]
  //: joint g22 (w39) @(234, 251) /w:[ 4 6 -1 3 ]
  //: joint g45 (w38) @(250, 510) /w:[ 16 18 -1 15 ]
  //: SWITCH g70 (w15) @(617,604) /sn:0 /w:[ 0 ] /st:0 /dn:0
  //: SWITCH g114 (w61) @(131,2131) /sn:0 /w:[ 1 ] /st:0 /dn:0
  H74182 g209 (._G0(w166), ._G1(w159), ._G2(w167), ._G3(w168), ._P0(w171), ._P1(w172), ._P2(w169), ._P3(w170), .Cn(w126), .CnPx(w164), .CnPy(w163), .CnPz(w162), ._G(w161), ._P(w160));   //: @(1090, 555) /sz:(105, 160) /sn:0 /p:[ Li0>1 Li1>0 Li2>1 Li3>0 Li4>1 Li5>1 Li6>1 Li7>0 Li8>1 Ro0<0 Ro1<0 Ro2<0 Ro3<0 Ro4<1 ]
  //: LED g229 (w177) @(426,1278) /sn:0 /w:[ 0 ] /type:0
  //: LED g30 (w22) @(459,183) /sn:0 /w:[ 0 ] /type:0
  //: joint g164 (w37) @(266, 990) /w:[ 26 25 -1 28 ]
  //: LED g118 (w103) @(886,1256) /sn:0 /w:[ 0 ] /type:0

endmodule
//: /netlistEnd

//: /hdlBegin H7442
//: interface  /sz:(89, 175) /bd:[ Li0>A0(16/175) Li1>A1(32/175) Li2>A2(48/175) Li3>A3(64/175) Ro0<_Y0(16/175) Ro1<_Y1(32/175) Ro2<_Y2(48/175) Ro3<_Y3(64/175) Ro4<_Y4(80/175) Ro5<_Y5(96/175) Ro6<_Y6(112/175) Ro7<_Y7(128/175) Ro8<_Y8(144/175) Ro9<_Y9(160/175) ] /pd: 0 /pi: 0 /pe: 1 /pp: 0
//: property pptype=0
//: enddecls
module H7442 #(.delay(14)) (A0,A1,A2,A3,_Y0,_Y1,_Y2,_Y3,_Y4,_Y5,_Y6,_Y7,_Y8,_Y9);
  input A0,A1,A2,A3;
  output _Y0,_Y1,_Y2,_Y3,_Y4,_Y5,_Y6,_Y7,_Y8,_Y9;
  wire c1_0, c1_1, c1_2, c1_3, c1_4, c1_5, c1_6;
  
  assign c1_0 = ~(~A0 & ~A1);
  assign c1_1 = ~(A0 & ~A1);
  assign c1_2 = ~(~A0 & A1);
  assign c1_3 = ~(A0 & A1);
  assign c1_4 = ~(~A2 & ~A3);
  assign c1_5 = ~(A2 & ~A3);
  assign c1_6 = ~(~A2 & A3);
  
  assign _Y0 = ~(~c1_0 & ~c1_4);
  assign _Y1 = ~(~c1_1 & ~c1_4);
  assign _Y2 = ~(~c1_2 & ~c1_4);
  assign _Y3 = ~(~c1_3 & ~c1_4);
  assign _Y4 = ~(~c1_0 & ~c1_5);
  assign _Y5 = ~(~c1_1 & ~c1_5);
  assign _Y6 = ~(~c1_2 & ~c1_5);
  assign _Y7 = ~(~c1_3 & ~c1_5);
  assign _Y8 = ~(~c1_0 & ~c1_6);
  assign _Y9 = ~(~c1_1 & ~c1_6);

endmodule
//: /hdlEnd


`timescale 1ns/1ns

//: /hdlBegin H74182
//: interface  /sz:(105, 160) /bd:[ Li0>Cn(144/160) Li1>_P3(128/160) Li2>_P2(112/160) Li3>_P1(96/160) Li4>_P0(80/160) Li5>_G3(64/160) Li6>_G2(48/160) Li7>_G1(32/160) Li8>_G0(16/160) Ro0<_P(80/160) Ro1<_G(64/160) Ro2<CnPz(48/160) Ro3<CnPy(32/160) Ro4<CnPx(16/160) ] /pd: 0 /pi: 0 /pe: 1 /pp: 0
//: property pptype=0
//: enddecls
module H74182 #(.delay(4)) (_G0,_G1,_G2,_G3,_P0,_P1,_P2,_P3,_P,_G,Cn,CnPx,CnPy,CnPz);
  
  input Cn;
  input _G0,_G1,_G2,_G3;
  input _P0,_P1,_P2,_P3;
  output _P,_G;
  output CnPx,CnPy,CnPz;
  
  assign #delay CnPx = ~( (_G0 & _P0) | (~Cn & _G0) );
  assign #delay CnPy = ~( (_G1 & _P1) | (_G0 & _G1 & _P0) | (~Cn & _G0 & _G1) );
  assign #delay CnPz = ~( (_G2 & _P2) | (_G1 & _G2 & _P1) | (_G0 & _G1 & _G2 & _P0) | (~Cn & _G0 & _G1 & _G2) );
  assign #delay _G = ~( (_G3 & _P3) | (_G2 & _G3 & _P2) | (_G1 & _G2 & _G3 & _P1) | ( _G0 & _G1 & _G2 & _G3) );
  assign #delay _P = _P0 | _P1 | _P2 | _P3; 

endmodule
//: /hdlEnd


`timescale 1ns/1ns

//: /hdlBegin H7474
//: interface  /sz:(110, 124) /bd:[ Li0>_CLR2(96/124) Li1>_PRE2(80/124) Li2>D2(64/124) Li3>_CLR1(48/124) Li4>_PRE1(32/124) Li5>D1(16/124) Bi0>CLK(54/110) Ro0<_Q2(64/124) Ro1<Q2(48/124) Ro2<_Q1(32/124) Ro3<Q1(16/124) ] /pd: 0 /pi: 0 /pe: 1 /pp: 0
//: property pptype=0
//: enddecls
module H7474 #(.delay(18)) (CLK,D1,_PRE1,_CLR1,D2,_PRE2,_CLR2,Q1,_Q1,Q2,_Q2);
  input CLK,D1,_PRE1,_CLR1,D2,_PRE2,_CLR2;
  output Q1,_Q1,Q2,_Q2;
  reg R1,R2;
  
  assign #delay _Q1 = ~R1;
  assign #delay _Q2 = ~R2;
  assign #delay Q1 = R1;
  assign #delay Q2 = R2;
  
  always @(negedge _PRE1 or negedge _CLR1)
    begin
      if (~_PRE1)
        R1 = 1'b1;
      else if (~_CLR1)
        R1 = 1'b0;
    end

  always @(negedge _PRE2 or negedge _CLR2)
    begin
      if (~_PRE2)
        R2 = 1'b1;
      else if (~_CLR2)
        R2 = 1'b0;
    end
  
  always @(posedge CLK)
    begin
      if (~_PRE1 && ~_CLR1)
        R1 = D1;
      if (~_PRE2 && ~_CLR2)
        R2 = D2;
    end
  
  
endmodule
//: /hdlEnd


`timescale 1ns/1ns

//: /hdlBegin H7404
//: interface  /sz:(74, 112) /bd:[ Li0>A6(96/112) Li1>A5(80/112) Li2>A4(64/112) Li3>A3(48/112) Li4>A2(32/112) Li5>A1(16/112) Ro0<Y6(96/112) Ro1<Y5(80/112) Ro2<Y4(64/112) Ro3<Y3(48/112) Ro4<Y2(32/112) Ro5<Y1(16/112) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
//: enddecls
module H7404 #(.delay(3)) (A1,A2,A3,A4,A5,A6,Y1,Y2,Y3,Y4,Y4,Y6);
  input A1,A2,A3,A4,A5,A6;
  output Y1,Y2,Y3,Y4,Y5,Y6;

  assign #delay Y1 = ~A1;
  assign #delay Y2 = ~A2;
  assign #delay Y3 = ~A3;
  assign #delay Y4 = ~A4;
  assign #delay Y5 = ~A5;
  assign #delay Y6 = ~A6;

endmodule
//: /hdlEnd


`timescale 1ns/1ns

//: /hdlBegin H7411
//: interface  /sz:(74, 160) /bd:[ Li0>A1(16/160) Li1>A2(32/160) Li2>A3(48/160) Li3>B1(64/160) Li4>B2(80/160) Li5>B3(96/160) Li6>C1(112/160) Li7>C2(128/160) Li8>C3(144/160) Ro0<Y1(16/160) Ro1<Y2(32/160) Ro2<Y3(48/160) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
//: enddecls
module H7411 #(.delay(6)) (A1,A2,A3,B1,B2,B3,C1,C2,C3,Y1,Y2,Y3);
  input A1,A2,A3,B1,B2,B3,C1,C2,C3;
  output Y1,Y2,Y3;
  
  assign #delay Y1 = A1 & B1 & C1;
  assign #delay Y2 = A2 & B2 & C2;
  assign #delay Y3 = A3 & B3 & C3;

endmodule
//: /hdlEnd


`timescale 1ns/1ns

//: /hdlBegin H7427
//: interface  /sz:(88, 160) /bd:[ Li0>A1(16/160) Li1>A2(32/160) Li2>A3(48/160) Li3>B1(64/160) Li4>B2(80/160) Li5>B3(96/160) Li6>C1(112/160) Li7>C2(128/160) Li8>C3(144/160) Ro0<Y1(16/160) Ro1<Y2(32/160) Ro2<Y3(48/160) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
//: enddecls
module H7427 #(.delay(6)) (A1,B1,C1,A2,B2,C2,A3,B3,C3,Y1,Y2,Y3);
  input A1,B1,C1,A2,B2,C2,A3,B3,C3;
  output Y1,Y2,Y3;
  
  assign #delay Y1 = ~(A1 | B1 | C1);
  assign #delay Y2 = ~(A2 | B2 | C2);
  assign #delay Y3 = ~(A3 | B3 | C3);
endmodule
//: /hdlEnd


`timescale 1ns/1ns

//: /hdlBegin H7420
//: interface  /sz:(74, 144) /bd:[ Li0>D2(128/144) Li1>D1(112/144) Li2>C2(96/144) Li3>C1(80/144) Li4>B2(64/144) Li5>B1(48/144) Li6>A2(32/144) Li7>A1(16/144) Ro0<Y2(32/144) Ro1<Y1(16/144) ] /pd: 0 /pi: 0 /pe: 0 /pp: 0
//: property pptype=0
//: enddecls
module H7420 #(.delay(6)) (A1,A2,B1,B2,C1,C2,D1,D2,Y1,Y2);
  input A1,A2,B1,B2,C1,C2,D1,D2;
  output Y1,Y2;
  
  assign #delay Y1 = ~(A1 & B1 & C1 & D1);
  assign #delay Y2 = ~(A2 & B2 & C2 & D2);

endmodule
//: /hdlEnd


`timescale 1ns/1ns

//: /hdlBegin H7402
//: interface  /sz:(74, 144) /bd:[ Li0>A1(16/144) Li1>A2(32/144) Li2>A3(48/144) Li3>A4(64/144) Li4>B1(80/144) Li5>B2(96/144) Li6>B3(112/144) Li7>B4(128/144) Ro0<Y1(16/144) Ro1<Y2(32/144) Ro2<Y3(48/144) Ro3<Y4(64/144) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
//: enddecls
module H7402 #(.delay(4)) (A1,A2,A3,A4,B1,B2,B3,B4,Y1,Y2,Y3,Y4);
  input A1,A2,A3,A4,B1,B2,B3,B4;
  output Y1,Y2,Y3,Y4;
  
  assign #delay Y1 = A1 ~| B1;
  assign #delay Y2 = A2 ~| B2;
  assign #delay Y3 = A3 ~| B3;
  assign #delay Y4 = A4 ~| B4;

endmodule
//: /hdlEnd


`timescale 1ns/1ns

//: /hdlBegin H74154
//: interface  /sz:(105, 272) /bd:[ Li0>_G2(96/272) Li1>_G1(80/272) Li2>D(64/272) Li3>C(48/272) Li4>B(32/272) Li5>A(16/272) Ro0<_Y16(256/272) Ro1<_Y15(240/272) Ro2<_Y14(224/272) Ro3<_Y13(208/272) Ro4<_Y12(192/272) Ro5<_Y11(176/272) Ro6<_Y10(160/272) Ro7<_Y9(144/272) Ro8<_Y8(128/272) Ro9<_Y7(112/272) Ro10<_Y6(96/272) Ro11<_Y5(80/272) Ro12<_Y4(64/272) Ro13<_Y3(48/272) Ro14<_Y2(32/272) Ro15<_Y1(16/272) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
//: enddecls
module H74154 #(.delay(20)) (A,B,C,D,_G1,_G2,_Y1,_Y2,_Y3,_Y4,_Y5,_Y6,_Y7,_Y8,
              _Y9,_Y10,_Y11,_Y12,_Y13,_Y14,_Y15,_Y16);
  input A,B,C,D,_G1,_G2;
  output _Y1,_Y2,_Y3,_Y4,_Y5,_Y6,_Y7,_Y8,_Y9,_Y10,_Y11,_Y12,_Y13,_Y14,_Y15,_Y16;
  reg [15:0] R;
  
  assign #delay {_Y16,_Y15,_Y14,_Y13,_Y12,_Y11,_Y10,_Y9,_Y8,_Y7,_Y6,_Y5,_Y4,_Y3,_Y2,_Y1} = ~R;

  initial
    if (_G1 || _G2)
      R = 0;
    else
      R = 16'h1 << {D,C,B,A};

  always @(_G1 or _G2 or A or B or C or D)
    if (_G1 || _G2)
      R = 0;
    else
      R = 16'h1 << {D,C,B,A};

endmodule
//: /hdlEnd


`timescale 1ns/1ns

//: /hdlBegin H74181
//: interface  /sz:(93, 240) /bd:[ Li0>S3(224/240) Li1>S2(208/240) Li2>S1(192/240) Li3>S0(176/240) Li4>M(160/240) Li5>Cn(144/240) Li6>_B3(128/240) Li7>_B2(112/240) Li8>_B1(96/240) Li9>_B0(80/240) Li10>_A3(64/240) Li11>_A2(48/240) Li12>_A1(32/240) Li13>_A0(16/240) Ro0<_P(128/240) Ro1<_G(112/240) Ro2<CnP4(96/240) Ro3<AEB(80/240) Ro4<_F3(64/240) Ro5<_F2(48/240) Ro6<_F1(32/240) Ro7<_F0(16/240) ] /pd: 0 /pi: 0 /pe: 1 /pp: 0
//: property pptype=0
//: enddecls
module H74181 #(.delay(4)) (_A0,_A1,_A2,_A3,_B0,_B1,_B2,_B3,S0,S1,S2,S3,Cn,M,_F0,_F1,_F2,_F3,AEB,CnP4,_G,_P);
  
  input _A0,_A1,_A2,_A3;
  input _B0,_B1,_B2,_B3;
  input Cn,M;
  input S0,S1,S2,S3;
  output _F0,_F1,_F2,_F3;
  output AEB,CnP4,_G,_P;
  
  // First level gates outputs
  wire L1_0,L1_1,L1_2,L1_3,L1_4,L1_5,L1_6,L1_7;
  
  assign #delay L1_0 = ~( _A0 | (_B0 & S0) | (~_B0 & S1) );
  assign #delay L1_1 = ~( (_A0 & ~_B0 & S2 ) | (_A0 & _B0 & S3) );
  
  assign #delay L1_2 = ~( _A1 | (_B1 & S0) | (~_B1 & S1) );
  assign #delay L1_3 = ~( (_A1 & ~_B1 & S2 ) | (_A1 & _B1 & S3) );
  
  assign #delay L1_4 = ~( _A2 | (_B2 & S0) | (~_B2 & S1) );
  assign #delay L1_5 = ~( (_A2 & ~_B2 & S2 ) | (_A2 & _B2 & S3) );
  
  assign #delay L1_6 = ~( _A3 | (_B3 & S0) | (~_B3 & S1) );
  assign #delay L1_7 = ~( (_A3 & ~_B3 & S2 ) | (_A3 & _B3 & S3) );
  
  // Second level gates output
  wire L2_0,L2_1,L2_2,L2_3;
  
  assign #delay L2_0 = ~(~M & Cn);
  assign #delay L2_1 = ~( (~M & L1_0) | (~M & L1_1 & Cn) );
  assign #delay L2_2 = ~( (~M & L1_2) | (~M & L1_0 & L1_3) | (~M & L1_1 & L1_3 & Cn)  );
  assign #delay L2_3 = ~( (~M & L1_4) | (~M & L1_2 & L1_5) | (~M & L1_0 & L1_3 & L1_5) | (~M & L1_1 & L1_3 & L1_5 &Cn)  );
  
  assign #delay _F0 = L2_0 ^ (L1_0 ^ L1_1);
  assign #delay _F1 = L2_1 ^ (L1_2 ^ L1_3); 
  assign #delay _F2 = L2_2 ^ (L1_4 ^ L1_5);
  assign #delay _F3 = L2_3 ^ (L1_6 ^ L1_7);
  
  assign #delay AEB = _F0 & _F1 & _F2 & _F3;
  assign #delay _G = ~( L1_6 | (L1_4 & L1_7) | (L1_2 & L1_5 & L1_7) | (L1_0 & L1_3 & L1_5 & L1_7) );
  assign #delay CnP4 = ~_G | ( L1_1 & L1_3 & L1_5 & L1_7 & Cn );
  assign #delay _P = ~( L1_1 & L1_3 & L1_5 & L1_7 );
    
endmodule
//: /hdlEnd


`timescale 1ns/1ns

//: /hdlBegin H74157
//: interface  /sz:(81, 176) /bd:[ Li0>S(160/176) Li1>_G(144/176) Li2>B4(128/176) Li3>B3(112/176) Li4>B2(96/176) Li5>B1(80/176) Li6>A4(64/176) Li7>A3(48/176) Li8>A2(32/176) Li9>A1(16/176) Ro0<Y4(64/176) Ro1<Y3(48/176) Ro2<Y2(32/176) Ro3<Y1(16/176) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
//: enddecls
module H74157 #(.delay(18)) (S,_G,A1,A2,A3,A4,B1,B2,B3,B4,Y1,Y2,Y3,Y4);
  input S,_G;
  input A1,A2,A3,A4,B1,B2,B3,B4;
  output Y1,Y2,Y3,Y4;
  
  assign #delay Y1 = _G ? 1'b1 : (S ? B1 : A1);
  assign #delay Y2 = _G ? 1'b1 : (S ? B2 : A2);
  assign #delay Y3 = _G ? 1'b1 : (S ? B3 : A3);
  assign #delay Y4 = _G ? 1'b1 : (S ? B4 : A4);

endmodule
//: /hdlEnd


`timescale 1ns/1ns

//: /hdlBegin H7486
//: interface  /sz:(74, 144) /bd:[ Li0>B4(128/144) Li1>B3(112/144) Li2>B2(96/144) Li3>B1(80/144) Li4>A4(64/144) Li5>A3(48/144) Li6>A2(32/144) Li7>A1(16/144) Ro0<Y4(64/144) Ro1<Y3(48/144) Ro2<Y2(32/144) Ro3<Y1(16/144) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
//: enddecls
module H7486 #(.delay(4)) (A1,A2,A3,A4,B1,B2,B3,B4,Y1,Y2,Y3,Y4);
  input A1,A2,A3,A4,B1,B2,B3,B4;
  output Y1,Y2,Y3,Y4;
  
  assign #delay Y1 = A1 ^ B1;
  assign #delay Y2 = A2 ^ B2;
  assign #delay Y3 = A3 ^ B3;
  assign #delay Y4 = A4 ^ B4;

endmodule
//: /hdlEnd


`timescale 1ns/1ns

//: /hdlBegin H7408
//: interface  /sz:(74, 144) /bd:[ Li0>A1(16/144) Li1>A2(32/144) Li2>A3(48/144) Li3>A4(64/144) Li4>B1(80/144) Li5>B2(96/144) Li6>B3(112/144) Li7>B4(128/144) Ro0<Y1(16/144) Ro1<Y2(32/144) Ro2<Y3(48/144) Ro3<Y4(64/144) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
//: enddecls
module H7408 #(.delay(4)) (A1,A2,A3,A4,B1,B2,B3,B4,Y1,Y2,Y3,Y4);
  input A1,A2,A3,A4,B1,B2,B3,B4;
  output Y1,Y2,Y3,Y4;
  
  assign #delay Y1 = A1 & B1;
  assign #delay Y2 = A2 & B2;
  assign #delay Y3 = A3 & B3;
  assign #delay Y4 = A4 & B4;

endmodule
//: /hdlEnd


`timescale 1ns/1ns

//: /hdlBegin H74163
//: interface  /sz:(117, 160) /bd:[ Li0>A(16/160) Li1>B(32/160) Li2>C(48/160) Li3>D(64/160) Li4>_CLR(80/160) Li5>ENP(96/160) Li6>ENT(112/160) Li7>_LOAD(128/160) Bi0>CLK(61/117) Ro0<QA(16/160) Ro1<QB(32/160) Ro2<QC(48/160) Ro3<QD(64/160) Ro4<RCO(80/160) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
//: enddecls
module H74163 #(.delay(20)) (_CLR, _LOAD, ENT, ENP, CLK, A, B, C, D, QA, QB, QC, QD, RCO);
  input _CLR, _LOAD, ENT, ENP, CLK, A, B, C, D;
  reg output QA, QB, QC, QD;
  output RCO;
  
  assign RCO = QA & QB & QC &QD & ENT;
  
  always @(_CLR or _LOAD)
    if (_CLR == 1'b0)
      begin
        QA <= #delay 1'b0;
        QB <= #delay 1'b0;
        QC <= #delay 1'b0;
        QD <= #delay 1'b0;
      end
    else if (_LOAD == 1'b0)
      begin
        QA <= #delay A;
        QB <= #delay B;
        QC <= #delay C;
        QD <= #delay D;
      end
  
  always @(posedge CLK)
    if (ENP == 1'b1 && ENT == 1'b1 && _CLR == 1'b1 && _LOAD == 1'b1)
      begin
        {QD, QC, QB, QA} <= #delay {QD, QC, QB, QA} + 4'h1;
      end

endmodule
//: /hdlEnd


`timescale 1ns/1ns

//: /hdlBegin H7410
//: interface  /sz:(74, 160) /bd:[ Li0>A1(16/160) Li1>A2(32/160) Li2>A3(48/160) Li3>B1(64/160) Li4>B2(80/160) Li5>B3(96/160) Li6>C1(112/160) Li7>C2(128/160) Li8>C3(144/160) Ro0<Y1(16/160) Ro1<Y2(32/160) Ro2<Y3(48/160) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
//: enddecls
module H7410 #(.delay(6)) (A1,A2,A3,B1,B2,B3,C1,C2,C3,Y1,Y2,Y3);
  input A1,A2,A3,B1,B2,B3,C1,C2,C3;
  output Y1,Y2,Y3;
  
  assign #delay Y1 = ~(A1 & B1 & C1);
  assign #delay Y2 = ~(A2 & B2 & C2);
  assign #delay Y3 = ~(A3 & B3 & C3);

endmodule
//: /hdlEnd


`timescale 1ns/1ns

//: /hdlBegin H74175
//: interface  /sz:(105, 144) /bd:[ Li0>D1(16/144) Li1>D2(32/144) Li2>D3(48/144) Li3>D4(64/144) Li4>_PRE(80/144) Li5>_CLR(96/144) Bi0>CLK(52/105) Ro0<Q1(16/144) Ro1<Q2(32/144) Ro2<Q3(48/144) Ro3<Q4(64/144) Ro4<_Q1(80/144) Ro5<_Q2(96/144) Ro6<_Q3(112/144) Ro7<_Q4(128/144) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
//: enddecls
module H74175 #(.delay(18)) (CLK,_PRE,_CLR,D1,D2,D3,D4,Q1,_Q1,Q2,_Q2,Q3,_Q3,Q4,_Q4);
  input CLK,_PRE,_CLR,D1,D2,D3,D4;
  output Q1,_Q1,Q2,_Q2,Q3,_Q3,Q4,_Q4;
  reg R1,R2,R3,R4;
  
  assign #delay _Q1 = ~R1;
  assign #delay _Q2 = ~R2;
  assign #delay _Q3 = ~R3;
  assign #delay _Q4 = ~R4;
  assign #delay Q1 = R1;
  assign #delay Q2 = R2;
  assign #delay Q3 = R3;
  assign #delay Q4 = R4;
  
  always @(negedge _PRE or negedge _CLR)
    begin
      if (~_PRE)
        begin
          R1 = 1'b1;
          R2 = 1'b1;
          R3 = 1'b1;
          R4 = 1'b1;
        end
      else if (~_CLR)
        begin
          R1 = 1'b0;
          R2 = 1'b0;
          R3 = 1'b0;
          R4 = 1'b0;
        end
    end

  always @(posedge CLK)
    begin
      if (~_PRE && ~_CLR)
        begin
          R1 = D1;
          R2 = D2;
          R3 = D3;
          R4 = D4;
        end
    end
  
  
endmodule
//: /hdlEnd


`timescale 1ns/1ns

//: /hdlBegin H7421
//: interface  /sz:(74, 144) /bd:[ Li0>D2(128/144) Li1>D1(112/144) Li2>C2(96/144) Li3>C1(80/144) Li4>B2(64/144) Li5>B1(48/144) Li6>A2(32/144) Li7>A1(16/144) Ro0<Y2(32/144) Ro1<Y1(16/144) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
//: enddecls
module H7421 #(.delay(6)) (A1,A2,B1,B2,C1,C2,D1,D2,Y1,Y2);
  input A1,A2,B1,B2,C1,C2,D1,D2;
  output Y1,Y2;
  
  assign #delay Y1 = A1 & B1 & C1 & D1;
  assign #delay Y2 = A2 & B2 & C2 & D2;

endmodule
//: /hdlEnd


`timescale 1ns/1ns

//: /hdlBegin H7430
//: interface  /sz:(62, 144) /bd:[ Li0>A(16/144) Li1>B(32/144) Li2>C(48/144) Li3>D(64/144) Li4>E(80/144) Li5>F(96/144) Li6>G(112/144) Li7>H(128/144) Ro0<Y(16/144) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
//: enddecls
module H7430 #(.delay(12)) (A,B,C,D,E,F,G,H,Y);
  input A,B,C,D,E,F,G,H;
  output Y;
  
  assign #delay Y = ~(A & B & C & D & E & F & G & H); 

endmodule
//: /hdlEnd


`timescale 1ns/1ns

//: /hdlBegin H7400
//: interface  /sz:(74, 144) /bd:[ Li0>A1(16/144) Li1>A2(32/144) Li2>A3(48/144) Li3>A4(64/144) Li4>B1(80/144) Li5>B2(96/144) Li6>B3(112/144) Li7>B4(128/144) Ro0<Y1(16/144) Ro1<Y2(32/144) Ro2<Y3(48/144) Ro3<Y4(64/144) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
//: enddecls
module H7400 #(.delay(4)) (A1,A2,A3,A4,B1,B2,B3,B4,Y1,Y2,Y3,Y4);
  input A1,A2,A3,A4,B1,B2,B3,B4;
  output Y1,Y2,Y3,Y4;
  
  assign #delay Y1 = A1 ~& B1;
  assign #delay Y2 = A2 ~& B2;
  assign #delay Y3 = A3 ~& B3;
  assign #delay Y4 = A4 ~& B4;

endmodule
//: /hdlEnd


`timescale 1ns/1ns

//: /hdlBegin H7432
//: interface  /sz:(74, 144) /bd:[ Li0>B4(128/144) Li1>B3(112/144) Li2>B2(96/144) Li3>B1(80/144) Li4>A4(64/144) Li5>A3(48/144) Li6>A2(32/144) Li7>A1(16/144) Ro0<Y4(64/144) Ro1<Y3(48/144) Ro2<Y2(32/144) Ro3<Y1(16/144) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
//: enddecls
module H7432 #(.delay(6)) (A1,A2,A3,A4,B1,B2,B3,B4,Y1,Y2,Y3,Y4);
  input A1,A2,A3,A4,B1,B2,B3,B4;
  output Y1,Y2,Y3,Y4;
  
  assign #delay Y1 = A1 | B1;
  assign #delay Y2 = A2 | B2;
  assign #delay Y3 = A3 | B3;
  assign #delay Y4 = A4 | B4;

endmodule
//: /hdlEnd


`timescale 1ns/1ns


//: version "2.2"
//: property encoding = "utf-8"
//: property locale = "uk"
//: property prefix = "_GG"
//: property title = "Сторінка підручника"
//: property showSwitchNets = 0
//: property discardChanges = 1
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin PAGE1
module PAGE1;    //: root_module
//: enddecls

  //: comment g1 @(475,291) /sn:0 /R:14 /anc:1
  //: /line:"<a href=\"welcome.v\">Повернутися до основної сторінки TkGate.</a>"
  //: /end
  //: comment g0 @(476,49) /sn:0 /anc:1
  //: /line:"<a href=\"welcome.v\"><img src=\"biggatelogo.gif\"></a>"
  //: /end
  //: comment g18 @(10,10) /sn:0 /anc:1
  //: /line:"<h1>Tutorial Chapters:</h1>"
  //: /line:""
  //: /line:"<h3><a href=\"create.v\">1. Створення схеми</a></h3> - Get started by creating a simple circuit."
  //: /line:""
  //: /line:"<h3><a href=\"gates.v\">2. Редагування шлюзів</a></h3> - The basics of editing gates."
  //: /line:""
  //: /line:"<h3><a href=\"wires.v\">3. Редагування дротів</a></h3> - The basics of editing wires."
  //: /line:""
  //: /line:"<h3><a href=\"group.v\">4. Можливості з редагування груп</a></h3> - Operate on groups of gates."
  //: /line:""
  //: /line:"<h3><a href=\"modules.v\">5. Використання модулів</a></h3> - Using modules in your circuit."
  //: /line:""
  //: /line:"<h3><a href=\"advanced.v\">6. Advanced Editing Techniques</a></h3> - Learn advanced editing tricks."
  //: /line:""
  //: /line:"<h3><a href=\"combinational1.v\">7. Комбінаційне моделювання</a></h3> - Simulate a circuit with"
  //: /line:"combinational logic."
  //: /line:""
  //: /line:"<h3><a href=\"sequential1.v\">8. Моделювання послідовності елементів</a></h3> - Simulate a circuit with sequential logic."
  //: /line:""
  //: /line:"<h3><a href=\"verilog.v\">9. Текстовий Verilog</a></h3> - Create modules with textual Verilog descriptions."
  //: /line:""
  //: /line:"<h3><a href=\"options.v\">10. Налаштовування TkGate</a></h3> - Customize TkGate to suit your tastes."
  //: /line:""
  //: /end

endmodule
//: /netlistEnd


//: version "2.1"
//: property encoding = "utf-8"
//: property locale = "ru"
//: property prefix = "_GG"
//: property title = "Настройка TkGate"
//: property showSwitchNets = 0
//: property discardChanges = 1
//: property timingViolationMode = 2
//: property initTime = "0 ns"
//: require "tty"

`timescale 1ns/1ns

//: /netlistBegin PAGE1
module PAGE1;    //: root_module
//: enddecls

  //: comment g1 @(219,134) /sn:0 /anc:1
  //: /line:"<img src=iface.gif>"
  //: /end
  //: comment g9 @(10,10) /anc:1
  //: /line:"<h3>Настройка TkGate</h3>"
  //: /line:""
  //: /line:"Этот раздел описывает некоторые настройки TkGate. Ваши настройки хранятся в файле"
  //: /line:"\".tkgate2-preferences\" в Вашем домашнем каталоге."
  //: /end
  //: comment g0 @(10,310) /sn:0 /anc:1
  //: /line:"<tutorial-navigation>"
  //: /end

endmodule
//: /netlistEnd

//: /netlistBegin PAGE3
module PAGE3();
//: interface  /sz:(40, 40) /bd:[ ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
//: enddecls

  //: comment g1 @(134,181) /sn:0 /anc:1
  //: /line:"<img src=example_bindings.gif>"
  //: /end
  //: comment g9 @(10,10) /anc:1
  //: /line:"<h3>Настройка TkGate</h3> <b>(изменение стиля назначения клавиш)</b>"
  //: /line:""
  //: /line:"Вы можете изменять стиль привязки клавиш в группе \"Интерфейс\" диалога настроек. В настоящее"
  //: /line:"время можно выбирать между стилями \"emacs\" и \"Windows\". Выбор стиля привязки сделает вызов"
  //: /line:"таких операций как копирование/вставка аналогичными Windows или Emacs. Однако, операции работы"
  //: /line:"с вентилями будут использовать одни и те же клавиши."
  //: /end
  //: comment g0 @(10,310) /sn:0
  //: /line:"<tutorial-navigation>"
  //: /end

endmodule
//: /netlistEnd

//: /netlistBegin PAGE2
module PAGE2();
//: interface  /sz:(40, 40) /bd:[ ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
//: enddecls

  //: comment g1 @(116,149) /sn:0 /anc:1
  //: /line:"<img src=example_name.gif>"
  //: /end
  //: comment g9 @(10,10) /anc:1
  //: /line:"<h3>Настрока TkGate</h3> <b>(Установка персональной идентификации)</b>"
  //: /line:""
  //: /line:"Для установки настроек TkGate, откройте диалог настроек, выбрав <font color=red2>Инструменты &rarr; Настройки</font> из меню. Введите имя компьютера"
  //: /line:"и Ваше собственное в разделе \"Общие\". Введённые значения будут использованы при печати из TkGate."
  //: /end
  //: comment g0 @(10,310) /sn:0 /anc:1
  //: /line:"<tutorial-navigation>"
  //: /end

endmodule
//: /netlistEnd


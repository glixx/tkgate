//: version "2.1-a2"
//: property encoding = "utf-8"
//: property locale = "de"
//: property prefix = "_GG"
//: property title = "sim_tut.v"
//: property useExtBars = 0
//: property discardChanges = 1

`timescale 1ns/1ns

//: /netlistBegin PAGE1
module PAGE1;    //: root_module
//: enddecls

  //: comment g13 @(10,10) /anc:1
  //: /line:"<h3>Simulation von Schaltnetzen</h3>"
  //: /line:""
  //: /line:"TkGate benutzt einen Verilog-basierten diskret-ereignisgesteuerten Simulator zur"
  //: /line:"Simulation der Schaltungsbeschreibung. In diesem Abschnitt werden die Grundlagen"
  //: /line:"beschrieben, die zur Simulation von Schaltnetzen benötigt werden."
  //: /end
  //: comment g0 @(191,165) /sn:0 /anc:1
  //: /line:"<img src=simulate.gif>"
  //: /end
  //: comment g12 @(10,410) /sn:0 /R:14 /anc:1
  //: /line:"<tutorial-navigation byfile=1>"
  //: /end

endmodule
//: /netlistEnd


`timescale 1ns/1ns

